module moji

// https://api.github.com/emojis

pub const db = map{
	':+1:': [byte(240),159,145,141]
	':-1:': [byte(240),159,145,142]
	':100:': [byte(240),159,146,175]
	':1234:': [byte(240),159,148,162]
	':1st_place_medal:': [byte(240),159,165,135]
	':2nd_place_medal:': [byte(240),159,165,136]
	':3rd_place_medal:': [byte(240),159,165,137]
	':8ball:': [byte(240),159,142,177]
	':a:': [byte(240),159,133,176]
	':ab:': [byte(240),159,134,142]
	':abacus:': [byte(240),159,167,174]
	':abc:': [byte(240),159,148,164]
	':abcd:': [byte(240),159,148,161]
	':accept:': [byte(240),159,137,145]
	':adhesive_bandage:': [byte(240),159,169,185]
	':adult:': [byte(240),159,167,145]
	':aerial_tramway:': [byte(240),159,154,161]
	':afghanistan:': [byte(240),159,135,166,240,159,135,171]
	':airplane:': [byte(226),156,136]
	':aland_islands:': [byte(240),159,135,166,240,159,135,189]
	':alarm_clock:': [byte(226),143,176]
	':albania:': [byte(240),159,135,166,240,159,135,177]
	':alembic:': [byte(226),154,151]
	':algeria:': [byte(240),159,135,169,240,159,135,191]
	':alien:': [byte(240),159,145,189]
	':ambulance:': [byte(240),159,154,145]
	':american_samoa:': [byte(240),159,135,166,240,159,135,184]
	':amphora:': [byte(240),159,143,186]
	':anchor:': [byte(226),154,147]
	':andorra:': [byte(240),159,135,166,240,159,135,169]
	':angel:': [byte(240),159,145,188]
	':anger:': [byte(240),159,146,162]
	':angola:': [byte(240),159,135,166,240,159,135,180]
	':angry:': [byte(240),159,152,160]
	':anguilla:': [byte(240),159,135,166,240,159,135,174]
	':anguished:': [byte(240),159,152,167]
	':ant:': [byte(240),159,144,156]
	':antarctica:': [byte(240),159,135,166,240,159,135,182]
	':antigua_barbuda:': [byte(240),159,135,166,240,159,135,172]
	':apple:': [byte(240),159,141,142]
	':aquarius:': [byte(226),153,146]
	':argentina:': [byte(240),159,135,166,240,159,135,183]
	':aries:': [byte(226),153,136]
	':armenia:': [byte(240),159,135,166,240,159,135,178]
	':arrow_backward:': [byte(226),151,128]
	':arrow_double_down:': [byte(226),143,172]
	':arrow_double_up:': [byte(226),143,171]
	':arrow_down:': [byte(226),172,135]
	':arrow_down_small:': [byte(240),159,148,189]
	':arrow_forward:': [byte(226),150,182]
	':arrow_heading_down:': [byte(226),164,181]
	':arrow_heading_up:': [byte(226),164,180]
	':arrow_left:': [byte(226),172,133]
	':arrow_lower_left:': [byte(226),134,153]
	':arrow_lower_right:': [byte(226),134,152]
	':arrow_right:': [byte(226),158,161]
	':arrow_right_hook:': [byte(226),134,170]
	':arrow_up:': [byte(226),172,134]
	':arrow_up_down:': [byte(226),134,149]
	':arrow_up_small:': [byte(240),159,148,188]
	':arrow_upper_left:': [byte(226),134,150]
	':arrow_upper_right:': [byte(226),134,151]
	':arrows_clockwise:': [byte(240),159,148,131]
	':arrows_counterclockwise:': [byte(240),159,148,132]
	':art:': [byte(240),159,142,168]
	':articulated_lorry:': [byte(240),159,154,155]
	':artificial_satellite:': [byte(240),159,155,176]
	':artist:': [byte(240),159,167,145,240,159,142,168]
	':aruba:': [byte(240),159,135,166,240,159,135,188]
	':ascension_island:': [byte(240),159,135,166,240,159,135,168]
	':asterisk:': [byte(42),226,131,163]
	':astonished:': [byte(240),159,152,178]
	':astronaut:': [byte(240),159,167,145,240,159,154,128]
	':athletic_shoe:': [byte(240),159,145,159]
	':atm:': [byte(240),159,143,167]
	':atom_symbol:': [byte(226),154,155]
	':australia:': [byte(240),159,135,166,240,159,135,186]
	':austria:': [byte(240),159,135,166,240,159,135,185]
	':auto_rickshaw:': [byte(240),159,155,186]
	':avocado:': [byte(240),159,165,145]
	':axe:': [byte(240),159,170,147]
	':azerbaijan:': [byte(240),159,135,166,240,159,135,191]
	':b:': [byte(240),159,133,177]
	':baby:': [byte(240),159,145,182]
	':baby_bottle:': [byte(240),159,141,188]
	':baby_chick:': [byte(240),159,144,164]
	':baby_symbol:': [byte(240),159,154,188]
	':back:': [byte(240),159,148,153]
	':bacon:': [byte(240),159,165,147]
	':badger:': [byte(240),159,166,161]
	':badminton:': [byte(240),159,143,184]
	':bagel:': [byte(240),159,165,175]
	':baggage_claim:': [byte(240),159,155,132]
	':baguette_bread:': [byte(240),159,165,150]
	':bahamas:': [byte(240),159,135,167,240,159,135,184]
	':bahrain:': [byte(240),159,135,167,240,159,135,173]
	':balance_scale:': [byte(226),154,150]
	':bald_man:': [byte(240),159,145,168,240,159,166,178]
	':bald_woman:': [byte(240),159,145,169,240,159,166,178]
	':ballet_shoes:': [byte(240),159,169,176]
	':balloon:': [byte(240),159,142,136]
	':ballot_box:': [byte(240),159,151,179]
	':ballot_box_with_check:': [byte(226),152,145]
	':bamboo:': [byte(240),159,142,141]
	':banana:': [byte(240),159,141,140]
	':bangbang:': [byte(226),128,188]
	':bangladesh:': [byte(240),159,135,167,240,159,135,169]
	':banjo:': [byte(240),159,170,149]
	':bank:': [byte(240),159,143,166]
	':bar_chart:': [byte(240),159,147,138]
	':barbados:': [byte(240),159,135,167,240,159,135,167]
	':barber:': [byte(240),159,146,136]
	':baseball:': [byte(226),154,190]
	':basket:': [byte(240),159,167,186]
	':basketball:': [byte(240),159,143,128]
	':basketball_man:': [byte(226),155,185,226,153,130]
	':basketball_woman:': [byte(226),155,185,226,153,128]
	':bat:': [byte(240),159,166,135]
	':bath:': [byte(240),159,155,128]
	':bathtub:': [byte(240),159,155,129]
	':battery:': [byte(240),159,148,139]
	':beach_umbrella:': [byte(240),159,143,150]
	':bear:': [byte(240),159,144,187]
	':bearded_person:': [byte(240),159,167,148]
	':bed:': [byte(240),159,155,143]
	':bee:': [byte(240),159,144,157]
	':beer:': [byte(240),159,141,186]
	':beers:': [byte(240),159,141,187]
	':beetle:': [byte(240),159,144,158]
	':beginner:': [byte(240),159,148,176]
	':belarus:': [byte(240),159,135,167,240,159,135,190]
	':belgium:': [byte(240),159,135,167,240,159,135,170]
	':belize:': [byte(240),159,135,167,240,159,135,191]
	':bell:': [byte(240),159,148,148]
	':bellhop_bell:': [byte(240),159,155,142]
	':benin:': [byte(240),159,135,167,240,159,135,175]
	':bento:': [byte(240),159,141,177]
	':bermuda:': [byte(240),159,135,167,240,159,135,178]
	':beverage_box:': [byte(240),159,167,131]
	':bhutan:': [byte(240),159,135,167,240,159,135,185]
	':bicyclist:': [byte(240),159,154,180]
	':bike:': [byte(240),159,154,178]
	':biking_man:': [byte(240),159,154,180,226,153,130]
	':biking_woman:': [byte(240),159,154,180,226,153,128]
	':bikini:': [byte(240),159,145,153]
	':billed_cap:': [byte(240),159,167,162]
	':biohazard:': [byte(226),152,163]
	':bird:': [byte(240),159,144,166]
	':birthday:': [byte(240),159,142,130]
	':black_circle:': [byte(226),154,171]
	':black_flag:': [byte(240),159,143,180]
	':black_heart:': [byte(240),159,150,164]
	':black_joker:': [byte(240),159,131,143]
	':black_large_square:': [byte(226),172,155]
	':black_medium_small_square:': [byte(226),151,190]
	':black_medium_square:': [byte(226),151,188]
	':black_nib:': [byte(226),156,146]
	':black_small_square:': [byte(226),150,170]
	':black_square_button:': [byte(240),159,148,178]
	':blond_haired_man:': [byte(240),159,145,177,226,153,130]
	':blond_haired_person:': [byte(240),159,145,177]
	':blond_haired_woman:': [byte(240),159,145,177,226,153,128]
	':blonde_woman:': [byte(240),159,145,177,226,153,128]
	':blossom:': [byte(240),159,140,188]
	':blowfish:': [byte(240),159,144,161]
	':blue_book:': [byte(240),159,147,152]
	':blue_car:': [byte(240),159,154,153]
	':blue_heart:': [byte(240),159,146,153]
	':blue_square:': [byte(240),159,159,166]
	':blush:': [byte(240),159,152,138]
	':boar:': [byte(240),159,144,151]
	':boat:': [byte(226),155,181]
	':bolivia:': [byte(240),159,135,167,240,159,135,180]
	':bomb:': [byte(240),159,146,163]
	':bone:': [byte(240),159,166,180]
	':book:': [byte(240),159,147,150]
	':bookmark:': [byte(240),159,148,150]
	':bookmark_tabs:': [byte(240),159,147,145]
	':books:': [byte(240),159,147,154]
	':boom:': [byte(240),159,146,165]
	':boot:': [byte(240),159,145,162]
	':bosnia_herzegovina:': [byte(240),159,135,167,240,159,135,166]
	':botswana:': [byte(240),159,135,167,240,159,135,188]
	':bouncing_ball_man:': [byte(226),155,185,226,153,130]
	':bouncing_ball_person:': [byte(226),155,185]
	':bouncing_ball_woman:': [byte(226),155,185,226,153,128]
	':bouquet:': [byte(240),159,146,144]
	':bouvet_island:': [byte(240),159,135,167,240,159,135,187]
	':bow:': [byte(240),159,153,135]
	':bow_and_arrow:': [byte(240),159,143,185]
	':bowing_man:': [byte(240),159,153,135,226,153,130]
	':bowing_woman:': [byte(240),159,153,135,226,153,128]
	':bowl_with_spoon:': [byte(240),159,165,163]
	':bowling:': [byte(240),159,142,179]
	':boxing_glove:': [byte(240),159,165,138]
	':boy:': [byte(240),159,145,166]
	':brain:': [byte(240),159,167,160]
	':brazil:': [byte(240),159,135,167,240,159,135,183]
	':bread:': [byte(240),159,141,158]
	':breast_feeding:': [byte(240),159,164,177]
	':bricks:': [byte(240),159,167,177]
	':bride_with_veil:': [byte(240),159,145,176]
	':bridge_at_night:': [byte(240),159,140,137]
	':briefcase:': [byte(240),159,146,188]
	':british_indian_ocean_territory:': [byte(240),159,135,174,240,159,135,180]
	':british_virgin_islands:': [byte(240),159,135,187,240,159,135,172]
	':broccoli:': [byte(240),159,165,166]
	':broken_heart:': [byte(240),159,146,148]
	':broom:': [byte(240),159,167,185]
	':brown_circle:': [byte(240),159,159,164]
	':brown_heart:': [byte(240),159,164,142]
	':brown_square:': [byte(240),159,159,171]
	':brunei:': [byte(240),159,135,167,240,159,135,179]
	':bug:': [byte(240),159,144,155]
	':building_construction:': [byte(240),159,143,151]
	':bulb:': [byte(240),159,146,161]
	':bulgaria:': [byte(240),159,135,167,240,159,135,172]
	':bullettrain_front:': [byte(240),159,154,133]
	':bullettrain_side:': [byte(240),159,154,132]
	':burkina_faso:': [byte(240),159,135,167,240,159,135,171]
	':burrito:': [byte(240),159,140,175]
	':burundi:': [byte(240),159,135,167,240,159,135,174]
	':bus:': [byte(240),159,154,140]
	':business_suit_levitating:': [byte(240),159,149,180]
	':busstop:': [byte(240),159,154,143]
	':bust_in_silhouette:': [byte(240),159,145,164]
	':busts_in_silhouette:': [byte(240),159,145,165]
	':butter:': [byte(240),159,167,136]
	':butterfly:': [byte(240),159,166,139]
	':cactus:': [byte(240),159,140,181]
	':cake:': [byte(240),159,141,176]
	':calendar:': [byte(240),159,147,134]
	':call_me_hand:': [byte(240),159,164,153]
	':calling:': [byte(240),159,147,178]
	':cambodia:': [byte(240),159,135,176,240,159,135,173]
	':camel:': [byte(240),159,144,171]
	':camera:': [byte(240),159,147,183]
	':camera_flash:': [byte(240),159,147,184]
	':cameroon:': [byte(240),159,135,168,240,159,135,178]
	':camping:': [byte(240),159,143,149]
	':canada:': [byte(240),159,135,168,240,159,135,166]
	':canary_islands:': [byte(240),159,135,174,240,159,135,168]
	':cancer:': [byte(226),153,139]
	':candle:': [byte(240),159,149,175]
	':candy:': [byte(240),159,141,172]
	':canned_food:': [byte(240),159,165,171]
	':canoe:': [byte(240),159,155,182]
	':cape_verde:': [byte(240),159,135,168,240,159,135,187]
	':capital_abcd:': [byte(240),159,148,160]
	':capricorn:': [byte(226),153,145]
	':car:': [byte(240),159,154,151]
	':card_file_box:': [byte(240),159,151,131]
	':card_index:': [byte(240),159,147,135]
	':card_index_dividers:': [byte(240),159,151,130]
	':caribbean_netherlands:': [byte(240),159,135,167,240,159,135,182]
	':carousel_horse:': [byte(240),159,142,160]
	':carrot:': [byte(240),159,165,149]
	':cartwheeling:': [byte(240),159,164,184]
	':cat:': [byte(240),159,144,177]
	':cat2:': [byte(240),159,144,136]
	':cayman_islands:': [byte(240),159,135,176,240,159,135,190]
	':cd:': [byte(240),159,146,191]
	':central_african_republic:': [byte(240),159,135,168,240,159,135,171]
	':ceuta_melilla:': [byte(240),159,135,170,240,159,135,166]
	':chad:': [byte(240),159,135,185,240,159,135,169]
	':chains:': [byte(226),155,147]
	':chair:': [byte(240),159,170,145]
	':champagne:': [byte(240),159,141,190]
	':chart:': [byte(240),159,146,185]
	':chart_with_downwards_trend:': [byte(240),159,147,137]
	':chart_with_upwards_trend:': [byte(240),159,147,136]
	':checkered_flag:': [byte(240),159,143,129]
	':cheese:': [byte(240),159,167,128]
	':cherries:': [byte(240),159,141,146]
	':cherry_blossom:': [byte(240),159,140,184]
	':chess_pawn:': [byte(226),153,159]
	':chestnut:': [byte(240),159,140,176]
	':chicken:': [byte(240),159,144,148]
	':child:': [byte(240),159,167,146]
	':children_crossing:': [byte(240),159,154,184]
	':chile:': [byte(240),159,135,168,240,159,135,177]
	':chipmunk:': [byte(240),159,144,191]
	':chocolate_bar:': [byte(240),159,141,171]
	':chopsticks:': [byte(240),159,165,162]
	':christmas_island:': [byte(240),159,135,168,240,159,135,189]
	':christmas_tree:': [byte(240),159,142,132]
	':church:': [byte(226),155,170]
	':cinema:': [byte(240),159,142,166]
	':circus_tent:': [byte(240),159,142,170]
	':city_sunrise:': [byte(240),159,140,135]
	':city_sunset:': [byte(240),159,140,134]
	':cityscape:': [byte(240),159,143,153]
	':cl:': [byte(240),159,134,145]
	':clamp:': [byte(240),159,151,156]
	':clap:': [byte(240),159,145,143]
	':clapper:': [byte(240),159,142,172]
	':classical_building:': [byte(240),159,143,155]
	':climbing:': [byte(240),159,167,151]
	':climbing_man:': [byte(240),159,167,151,226,153,130]
	':climbing_woman:': [byte(240),159,167,151,226,153,128]
	':clinking_glasses:': [byte(240),159,165,130]
	':clipboard:': [byte(240),159,147,139]
	':clipperton_island:': [byte(240),159,135,168,240,159,135,181]
	':clock1:': [byte(240),159,149,144]
	':clock10:': [byte(240),159,149,153]
	':clock1030:': [byte(240),159,149,165]
	':clock11:': [byte(240),159,149,154]
	':clock1130:': [byte(240),159,149,166]
	':clock12:': [byte(240),159,149,155]
	':clock1230:': [byte(240),159,149,167]
	':clock130:': [byte(240),159,149,156]
	':clock2:': [byte(240),159,149,145]
	':clock230:': [byte(240),159,149,157]
	':clock3:': [byte(240),159,149,146]
	':clock330:': [byte(240),159,149,158]
	':clock4:': [byte(240),159,149,147]
	':clock430:': [byte(240),159,149,159]
	':clock5:': [byte(240),159,149,148]
	':clock530:': [byte(240),159,149,160]
	':clock6:': [byte(240),159,149,149]
	':clock630:': [byte(240),159,149,161]
	':clock7:': [byte(240),159,149,150]
	':clock730:': [byte(240),159,149,162]
	':clock8:': [byte(240),159,149,151]
	':clock830:': [byte(240),159,149,163]
	':clock9:': [byte(240),159,149,152]
	':clock930:': [byte(240),159,149,164]
	':closed_book:': [byte(240),159,147,149]
	':closed_lock_with_key:': [byte(240),159,148,144]
	':closed_umbrella:': [byte(240),159,140,130]
	':cloud:': [byte(226),152,129]
	':cloud_with_lightning:': [byte(240),159,140,169]
	':cloud_with_lightning_and_rain:': [byte(226),155,136]
	':cloud_with_rain:': [byte(240),159,140,167]
	':cloud_with_snow:': [byte(240),159,140,168]
	':clown_face:': [byte(240),159,164,161]
	':clubs:': [byte(226),153,163]
	':cn:': [byte(240),159,135,168,240,159,135,179]
	':coat:': [byte(240),159,167,165]
	':cocktail:': [byte(240),159,141,184]
	':coconut:': [byte(240),159,165,165]
	':cocos_islands:': [byte(240),159,135,168,240,159,135,168]
	':coffee:': [byte(226),152,149]
	':coffin:': [byte(226),154,176]
	':cold_face:': [byte(240),159,165,182]
	':cold_sweat:': [byte(240),159,152,176]
	':collision:': [byte(240),159,146,165]
	':colombia:': [byte(240),159,135,168,240,159,135,180]
	':comet:': [byte(226),152,132]
	':comoros:': [byte(240),159,135,176,240,159,135,178]
	':compass:': [byte(240),159,167,173]
	':computer:': [byte(240),159,146,187]
	':computer_mouse:': [byte(240),159,150,177]
	':confetti_ball:': [byte(240),159,142,138]
	':confounded:': [byte(240),159,152,150]
	':confused:': [byte(240),159,152,149]
	':congo_brazzaville:': [byte(240),159,135,168,240,159,135,172]
	':congo_kinshasa:': [byte(240),159,135,168,240,159,135,169]
	':congratulations:': [byte(227),138,151]
	':construction:': [byte(240),159,154,167]
	':construction_worker:': [byte(240),159,145,183]
	':construction_worker_man:': [byte(240),159,145,183,226,153,130]
	':construction_worker_woman:': [byte(240),159,145,183,226,153,128]
	':control_knobs:': [byte(240),159,142,155]
	':convenience_store:': [byte(240),159,143,170]
	':cook:': [byte(240),159,167,145,240,159,141,179]
	':cook_islands:': [byte(240),159,135,168,240,159,135,176]
	':cookie:': [byte(240),159,141,170]
	':cool:': [byte(240),159,134,146]
	':cop:': [byte(240),159,145,174]
	':copyright:': [byte(194),169]
	':corn:': [byte(240),159,140,189]
	':costa_rica:': [byte(240),159,135,168,240,159,135,183]
	':cote_divoire:': [byte(240),159,135,168,240,159,135,174]
	':couch_and_lamp:': [byte(240),159,155,139]
	':couple:': [byte(240),159,145,171]
	':couple_with_heart:': [byte(240),159,146,145]
	':couple_with_heart_man_man:': [byte(240),159,145,168,226,157,164,240,159,145,168]
	':couple_with_heart_woman_man:': [byte(240),159,145,169,226,157,164,240,159,145,168]
	':couple_with_heart_woman_woman:': [byte(240),159,145,169,226,157,164,240,159,145,169]
	':couplekiss:': [byte(240),159,146,143]
	':couplekiss_man_man:': [byte(240),159,145,168,226,157,164,240,159,146,139,240,159,145,168]
	':couplekiss_man_woman:': [byte(240),159,145,169,226,157,164,240,159,146,139,240,159,145,168]
	':couplekiss_woman_woman:': [byte(240),159,145,169,226,157,164,240,159,146,139,240,159,145,169]
	':cow:': [byte(240),159,144,174]
	':cow2:': [byte(240),159,144,132]
	':cowboy_hat_face:': [byte(240),159,164,160]
	':crab:': [byte(240),159,166,128]
	':crayon:': [byte(240),159,150,141]
	':credit_card:': [byte(240),159,146,179]
	':crescent_moon:': [byte(240),159,140,153]
	':cricket:': [byte(240),159,166,151]
	':cricket_game:': [byte(240),159,143,143]
	':croatia:': [byte(240),159,135,173,240,159,135,183]
	':crocodile:': [byte(240),159,144,138]
	':croissant:': [byte(240),159,165,144]
	':crossed_fingers:': [byte(240),159,164,158]
	':crossed_flags:': [byte(240),159,142,140]
	':crossed_swords:': [byte(226),154,148]
	':crown:': [byte(240),159,145,145]
	':cry:': [byte(240),159,152,162]
	':crying_cat_face:': [byte(240),159,152,191]
	':crystal_ball:': [byte(240),159,148,174]
	':cuba:': [byte(240),159,135,168,240,159,135,186]
	':cucumber:': [byte(240),159,165,146]
	':cup_with_straw:': [byte(240),159,165,164]
	':cupcake:': [byte(240),159,167,129]
	':cupid:': [byte(240),159,146,152]
	':curacao:': [byte(240),159,135,168,240,159,135,188]
	':curling_stone:': [byte(240),159,165,140]
	':curly_haired_man:': [byte(240),159,145,168,240,159,166,177]
	':curly_haired_woman:': [byte(240),159,145,169,240,159,166,177]
	':curly_loop:': [byte(226),158,176]
	':currency_exchange:': [byte(240),159,146,177]
	':curry:': [byte(240),159,141,155]
	':cursing_face:': [byte(240),159,164,172]
	':custard:': [byte(240),159,141,174]
	':customs:': [byte(240),159,155,131]
	':cut_of_meat:': [byte(240),159,165,169]
	':cyclone:': [byte(240),159,140,128]
	':cyprus:': [byte(240),159,135,168,240,159,135,190]
	':czech_republic:': [byte(240),159,135,168,240,159,135,191]
	':dagger:': [byte(240),159,151,161]
	':dancer:': [byte(240),159,146,131]
	':dancers:': [byte(240),159,145,175]
	':dancing_men:': [byte(240),159,145,175,226,153,130]
	':dancing_women:': [byte(240),159,145,175,226,153,128]
	':dango:': [byte(240),159,141,161]
	':dark_sunglasses:': [byte(240),159,149,182]
	':dart:': [byte(240),159,142,175]
	':dash:': [byte(240),159,146,168]
	':date:': [byte(240),159,147,133]
	':de:': [byte(240),159,135,169,240,159,135,170]
	':deaf_man:': [byte(240),159,167,143,226,153,130]
	':deaf_person:': [byte(240),159,167,143]
	':deaf_woman:': [byte(240),159,167,143,226,153,128]
	':deciduous_tree:': [byte(240),159,140,179]
	':deer:': [byte(240),159,166,140]
	':denmark:': [byte(240),159,135,169,240,159,135,176]
	':department_store:': [byte(240),159,143,172]
	':derelict_house:': [byte(240),159,143,154]
	':desert:': [byte(240),159,143,156]
	':desert_island:': [byte(240),159,143,157]
	':desktop_computer:': [byte(240),159,150,165]
	':detective:': [byte(240),159,149,181]
	':diamond_shape_with_a_dot_inside:': [byte(240),159,146,160]
	':diamonds:': [byte(226),153,166]
	':diego_garcia:': [byte(240),159,135,169,240,159,135,172]
	':disappointed:': [byte(240),159,152,158]
	':disappointed_relieved:': [byte(240),159,152,165]
	':diving_mask:': [byte(240),159,164,191]
	':diya_lamp:': [byte(240),159,170,148]
	':dizzy:': [byte(240),159,146,171]
	':dizzy_face:': [byte(240),159,152,181]
	':djibouti:': [byte(240),159,135,169,240,159,135,175]
	':dna:': [byte(240),159,167,172]
	':do_not_litter:': [byte(240),159,154,175]
	':dog:': [byte(240),159,144,182]
	':dog2:': [byte(240),159,144,149]
	':dollar:': [byte(240),159,146,181]
	':dolls:': [byte(240),159,142,142]
	':dolphin:': [byte(240),159,144,172]
	':dominica:': [byte(240),159,135,169,240,159,135,178]
	':dominican_republic:': [byte(240),159,135,169,240,159,135,180]
	':door:': [byte(240),159,154,170]
	':doughnut:': [byte(240),159,141,169]
	':dove:': [byte(240),159,149,138]
	':dragon:': [byte(240),159,144,137]
	':dragon_face:': [byte(240),159,144,178]
	':dress:': [byte(240),159,145,151]
	':dromedary_camel:': [byte(240),159,144,170]
	':drooling_face:': [byte(240),159,164,164]
	':drop_of_blood:': [byte(240),159,169,184]
	':droplet:': [byte(240),159,146,167]
	':drum:': [byte(240),159,165,129]
	':duck:': [byte(240),159,166,134]
	':dumpling:': [byte(240),159,165,159]
	':dvd:': [byte(240),159,147,128]
	':e-mail:': [byte(240),159,147,167]
	':eagle:': [byte(240),159,166,133]
	':ear:': [byte(240),159,145,130]
	':ear_of_rice:': [byte(240),159,140,190]
	':ear_with_hearing_aid:': [byte(240),159,166,187]
	':earth_africa:': [byte(240),159,140,141]
	':earth_americas:': [byte(240),159,140,142]
	':earth_asia:': [byte(240),159,140,143]
	':ecuador:': [byte(240),159,135,170,240,159,135,168]
	':egg:': [byte(240),159,165,154]
	':eggplant:': [byte(240),159,141,134]
	':egypt:': [byte(240),159,135,170,240,159,135,172]
	':eight:': [byte(56),226,131,163]
	':eight_pointed_black_star:': [byte(226),156,180]
	':eight_spoked_asterisk:': [byte(226),156,179]
	':eject_button:': [byte(226),143,143]
	':el_salvador:': [byte(240),159,135,184,240,159,135,187]
	':electric_plug:': [byte(240),159,148,140]
	':elephant:': [byte(240),159,144,152]
	':elf:': [byte(240),159,167,157]
	':elf_man:': [byte(240),159,167,157,226,153,130]
	':elf_woman:': [byte(240),159,167,157,226,153,128]
	':email:': [byte(226),156,137]
	':end:': [byte(240),159,148,154]
	':england:': [byte(240),159,143,180,243,160,129,167,243,160,129,162,243,160,129,165,243,160,129,174,243,160,129,167,243,160,129,191]
	':envelope:': [byte(226),156,137]
	':envelope_with_arrow:': [byte(240),159,147,169]
	':equatorial_guinea:': [byte(240),159,135,172,240,159,135,182]
	':eritrea:': [byte(240),159,135,170,240,159,135,183]
	':es:': [byte(240),159,135,170,240,159,135,184]
	':estonia:': [byte(240),159,135,170,240,159,135,170]
	':ethiopia:': [byte(240),159,135,170,240,159,135,185]
	':eu:': [byte(240),159,135,170,240,159,135,186]
	':euro:': [byte(240),159,146,182]
	':european_castle:': [byte(240),159,143,176]
	':european_post_office:': [byte(240),159,143,164]
	':european_union:': [byte(240),159,135,170,240,159,135,186]
	':evergreen_tree:': [byte(240),159,140,178]
	':exclamation:': [byte(226),157,151]
	':exploding_head:': [byte(240),159,164,175]
	':expressionless:': [byte(240),159,152,145]
	':eye:': [byte(240),159,145,129]
	':eye_speech_bubble:': [byte(240),159,145,129,240,159,151,168]
	':eyeglasses:': [byte(240),159,145,147]
	':eyes:': [byte(240),159,145,128]
	':face_with_head_bandage:': [byte(240),159,164,149]
	':face_with_thermometer:': [byte(240),159,164,146]
	':facepalm:': [byte(240),159,164,166]
	':facepunch:': [byte(240),159,145,138]
	':factory:': [byte(240),159,143,173]
	':factory_worker:': [byte(240),159,167,145,240,159,143,173]
	':fairy:': [byte(240),159,167,154]
	':fairy_man:': [byte(240),159,167,154,226,153,130]
	':fairy_woman:': [byte(240),159,167,154,226,153,128]
	':falafel:': [byte(240),159,167,134]
	':falkland_islands:': [byte(240),159,135,171,240,159,135,176]
	':fallen_leaf:': [byte(240),159,141,130]
	':family:': [byte(240),159,145,170]
	':family_man_boy:': [byte(240),159,145,168,240,159,145,166]
	':family_man_boy_boy:': [byte(240),159,145,168,240,159,145,166,240,159,145,166]
	':family_man_girl:': [byte(240),159,145,168,240,159,145,167]
	':family_man_girl_boy:': [byte(240),159,145,168,240,159,145,167,240,159,145,166]
	':family_man_girl_girl:': [byte(240),159,145,168,240,159,145,167,240,159,145,167]
	':family_man_man_boy:': [byte(240),159,145,168,240,159,145,168,240,159,145,166]
	':family_man_man_boy_boy:': [byte(240),159,145,168,240,159,145,168,240,159,145,166,240,159,145,166]
	':family_man_man_girl:': [byte(240),159,145,168,240,159,145,168,240,159,145,167]
	':family_man_man_girl_boy:': [byte(240),159,145,168,240,159,145,168,240,159,145,167,240,159,145,166]
	':family_man_man_girl_girl:': [byte(240),159,145,168,240,159,145,168,240,159,145,167,240,159,145,167]
	':family_man_woman_boy:': [byte(240),159,145,168,240,159,145,169,240,159,145,166]
	':family_man_woman_boy_boy:': [byte(240),159,145,168,240,159,145,169,240,159,145,166,240,159,145,166]
	':family_man_woman_girl:': [byte(240),159,145,168,240,159,145,169,240,159,145,167]
	':family_man_woman_girl_boy:': [byte(240),159,145,168,240,159,145,169,240,159,145,167,240,159,145,166]
	':family_man_woman_girl_girl:': [byte(240),159,145,168,240,159,145,169,240,159,145,167,240,159,145,167]
	':family_woman_boy:': [byte(240),159,145,169,240,159,145,166]
	':family_woman_boy_boy:': [byte(240),159,145,169,240,159,145,166,240,159,145,166]
	':family_woman_girl:': [byte(240),159,145,169,240,159,145,167]
	':family_woman_girl_boy:': [byte(240),159,145,169,240,159,145,167,240,159,145,166]
	':family_woman_girl_girl:': [byte(240),159,145,169,240,159,145,167,240,159,145,167]
	':family_woman_woman_boy:': [byte(240),159,145,169,240,159,145,169,240,159,145,166]
	':family_woman_woman_boy_boy:': [byte(240),159,145,169,240,159,145,169,240,159,145,166,240,159,145,166]
	':family_woman_woman_girl:': [byte(240),159,145,169,240,159,145,169,240,159,145,167]
	':family_woman_woman_girl_boy:': [byte(240),159,145,169,240,159,145,169,240,159,145,167,240,159,145,166]
	':family_woman_woman_girl_girl:': [byte(240),159,145,169,240,159,145,169,240,159,145,167,240,159,145,167]
	':farmer:': [byte(240),159,167,145,240,159,140,190]
	':faroe_islands:': [byte(240),159,135,171,240,159,135,180]
	':fast_forward:': [byte(226),143,169]
	':fax:': [byte(240),159,147,160]
	':fearful:': [byte(240),159,152,168]
	':feet:': [byte(240),159,144,190]
	':female_detective:': [byte(240),159,149,181,226,153,128]
	':female_sign:': [byte(226),153,128]
	':ferris_wheel:': [byte(240),159,142,161]
	':ferry:': [byte(226),155,180]
	':field_hockey:': [byte(240),159,143,145]
	':fiji:': [byte(240),159,135,171,240,159,135,175]
	':file_cabinet:': [byte(240),159,151,132]
	':file_folder:': [byte(240),159,147,129]
	':film_projector:': [byte(240),159,147,189]
	':film_strip:': [byte(240),159,142,158]
	':finland:': [byte(240),159,135,171,240,159,135,174]
	':fire:': [byte(240),159,148,165]
	':fire_engine:': [byte(240),159,154,146]
	':fire_extinguisher:': [byte(240),159,167,175]
	':firecracker:': [byte(240),159,167,168]
	':firefighter:': [byte(240),159,167,145,240,159,154,146]
	':fireworks:': [byte(240),159,142,134]
	':first_quarter_moon:': [byte(240),159,140,147]
	':first_quarter_moon_with_face:': [byte(240),159,140,155]
	':fish:': [byte(240),159,144,159]
	':fish_cake:': [byte(240),159,141,165]
	':fishing_pole_and_fish:': [byte(240),159,142,163]
	':fist:': [byte(226),156,138]
	':fist_left:': [byte(240),159,164,155]
	':fist_oncoming:': [byte(240),159,145,138]
	':fist_raised:': [byte(226),156,138]
	':fist_right:': [byte(240),159,164,156]
	':five:': [byte(53),226,131,163]
	':flags:': [byte(240),159,142,143]
	':flamingo:': [byte(240),159,166,169]
	':flashlight:': [byte(240),159,148,166]
	':flat_shoe:': [byte(240),159,165,191]
	':fleur_de_lis:': [byte(226),154,156]
	':flight_arrival:': [byte(240),159,155,172]
	':flight_departure:': [byte(240),159,155,171]
	':flipper:': [byte(240),159,144,172]
	':floppy_disk:': [byte(240),159,146,190]
	':flower_playing_cards:': [byte(240),159,142,180]
	':flushed:': [byte(240),159,152,179]
	':flying_disc:': [byte(240),159,165,143]
	':flying_saucer:': [byte(240),159,155,184]
	':fog:': [byte(240),159,140,171]
	':foggy:': [byte(240),159,140,129]
	':foot:': [byte(240),159,166,182]
	':football:': [byte(240),159,143,136]
	':footprints:': [byte(240),159,145,163]
	':fork_and_knife:': [byte(240),159,141,180]
	':fortune_cookie:': [byte(240),159,165,160]
	':fountain:': [byte(226),155,178]
	':fountain_pen:': [byte(240),159,150,139]
	':four:': [byte(52),226,131,163]
	':four_leaf_clover:': [byte(240),159,141,128]
	':fox_face:': [byte(240),159,166,138]
	':fr:': [byte(240),159,135,171,240,159,135,183]
	':framed_picture:': [byte(240),159,150,188]
	':free:': [byte(240),159,134,147]
	':french_guiana:': [byte(240),159,135,172,240,159,135,171]
	':french_polynesia:': [byte(240),159,135,181,240,159,135,171]
	':french_southern_territories:': [byte(240),159,135,185,240,159,135,171]
	':fried_egg:': [byte(240),159,141,179]
	':fried_shrimp:': [byte(240),159,141,164]
	':fries:': [byte(240),159,141,159]
	':frog:': [byte(240),159,144,184]
	':frowning:': [byte(240),159,152,166]
	':frowning_face:': [byte(226),152,185]
	':frowning_man:': [byte(240),159,153,141,226,153,130]
	':frowning_person:': [byte(240),159,153,141]
	':frowning_woman:': [byte(240),159,153,141,226,153,128]
	':fu:': [byte(240),159,150,149]
	':fuelpump:': [byte(226),155,189]
	':full_moon:': [byte(240),159,140,149]
	':full_moon_with_face:': [byte(240),159,140,157]
	':funeral_urn:': [byte(226),154,177]
	':gabon:': [byte(240),159,135,172,240,159,135,166]
	':gambia:': [byte(240),159,135,172,240,159,135,178]
	':game_die:': [byte(240),159,142,178]
	':garlic:': [byte(240),159,167,132]
	':gb:': [byte(240),159,135,172,240,159,135,167]
	':gear:': [byte(226),154,153]
	':gem:': [byte(240),159,146,142]
	':gemini:': [byte(226),153,138]
	':genie:': [byte(240),159,167,158]
	':genie_man:': [byte(240),159,167,158,226,153,130]
	':genie_woman:': [byte(240),159,167,158,226,153,128]
	':georgia:': [byte(240),159,135,172,240,159,135,170]
	':ghana:': [byte(240),159,135,172,240,159,135,173]
	':ghost:': [byte(240),159,145,187]
	':gibraltar:': [byte(240),159,135,172,240,159,135,174]
	':gift:': [byte(240),159,142,129]
	':gift_heart:': [byte(240),159,146,157]
	':giraffe:': [byte(240),159,166,146]
	':girl:': [byte(240),159,145,167]
	':globe_with_meridians:': [byte(240),159,140,144]
	':gloves:': [byte(240),159,167,164]
	':goal_net:': [byte(240),159,165,133]
	':goat:': [byte(240),159,144,144]
	':goggles:': [byte(240),159,165,189]
	':golf:': [byte(226),155,179]
	':golfing:': [byte(240),159,143,140]
	':golfing_man:': [byte(240),159,143,140,226,153,130]
	':golfing_woman:': [byte(240),159,143,140,226,153,128]
	':gorilla:': [byte(240),159,166,141]
	':grapes:': [byte(240),159,141,135]
	':greece:': [byte(240),159,135,172,240,159,135,183]
	':green_apple:': [byte(240),159,141,143]
	':green_book:': [byte(240),159,147,151]
	':green_circle:': [byte(240),159,159,162]
	':green_heart:': [byte(240),159,146,154]
	':green_salad:': [byte(240),159,165,151]
	':green_square:': [byte(240),159,159,169]
	':greenland:': [byte(240),159,135,172,240,159,135,177]
	':grenada:': [byte(240),159,135,172,240,159,135,169]
	':grey_exclamation:': [byte(226),157,149]
	':grey_question:': [byte(226),157,148]
	':grimacing:': [byte(240),159,152,172]
	':grin:': [byte(240),159,152,129]
	':grinning:': [byte(240),159,152,128]
	':guadeloupe:': [byte(240),159,135,172,240,159,135,181]
	':guam:': [byte(240),159,135,172,240,159,135,186]
	':guard:': [byte(240),159,146,130]
	':guardsman:': [byte(240),159,146,130,226,153,130]
	':guardswoman:': [byte(240),159,146,130,226,153,128]
	':guatemala:': [byte(240),159,135,172,240,159,135,185]
	':guernsey:': [byte(240),159,135,172,240,159,135,172]
	':guide_dog:': [byte(240),159,166,174]
	':guinea:': [byte(240),159,135,172,240,159,135,179]
	':guinea_bissau:': [byte(240),159,135,172,240,159,135,188]
	':guitar:': [byte(240),159,142,184]
	':gun:': [byte(240),159,148,171]
	':guyana:': [byte(240),159,135,172,240,159,135,190]
	':haircut:': [byte(240),159,146,135]
	':haircut_man:': [byte(240),159,146,135,226,153,130]
	':haircut_woman:': [byte(240),159,146,135,226,153,128]
	':haiti:': [byte(240),159,135,173,240,159,135,185]
	':hamburger:': [byte(240),159,141,148]
	':hammer:': [byte(240),159,148,168]
	':hammer_and_pick:': [byte(226),154,146]
	':hammer_and_wrench:': [byte(240),159,155,160]
	':hamster:': [byte(240),159,144,185]
	':hand:': [byte(226),156,139]
	':hand_over_mouth:': [byte(240),159,164,173]
	':handbag:': [byte(240),159,145,156]
	':handball_person:': [byte(240),159,164,190]
	':handshake:': [byte(240),159,164,157]
	':hankey:': [byte(240),159,146,169]
	':hash:': [byte(35),226,131,163]
	':hatched_chick:': [byte(240),159,144,165]
	':hatching_chick:': [byte(240),159,144,163]
	':headphones:': [byte(240),159,142,167]
	':health_worker:': [byte(240),159,167,145,226,154,149]
	':hear_no_evil:': [byte(240),159,153,137]
	':heard_mcdonald_islands:': [byte(240),159,135,173,240,159,135,178]
	':heart:': [byte(226),157,164]
	':heart_decoration:': [byte(240),159,146,159]
	':heart_eyes:': [byte(240),159,152,141]
	':heart_eyes_cat:': [byte(240),159,152,187]
	':heartbeat:': [byte(240),159,146,147]
	':heartpulse:': [byte(240),159,146,151]
	':hearts:': [byte(226),153,165]
	':heavy_check_mark:': [byte(226),156,148]
	':heavy_division_sign:': [byte(226),158,151]
	':heavy_dollar_sign:': [byte(240),159,146,178]
	':heavy_exclamation_mark:': [byte(226),157,151]
	':heavy_heart_exclamation:': [byte(226),157,163]
	':heavy_minus_sign:': [byte(226),158,150]
	':heavy_multiplication_x:': [byte(226),156,150]
	':heavy_plus_sign:': [byte(226),158,149]
	':hedgehog:': [byte(240),159,166,148]
	':helicopter:': [byte(240),159,154,129]
	':herb:': [byte(240),159,140,191]
	':hibiscus:': [byte(240),159,140,186]
	':high_brightness:': [byte(240),159,148,134]
	':high_heel:': [byte(240),159,145,160]
	':hiking_boot:': [byte(240),159,165,190]
	':hindu_temple:': [byte(240),159,155,149]
	':hippopotamus:': [byte(240),159,166,155]
	':hocho:': [byte(240),159,148,170]
	':hole:': [byte(240),159,149,179]
	':honduras:': [byte(240),159,135,173,240,159,135,179]
	':honey_pot:': [byte(240),159,141,175]
	':honeybee:': [byte(240),159,144,157]
	':hong_kong:': [byte(240),159,135,173,240,159,135,176]
	':horse:': [byte(240),159,144,180]
	':horse_racing:': [byte(240),159,143,135]
	':hospital:': [byte(240),159,143,165]
	':hot_face:': [byte(240),159,165,181]
	':hot_pepper:': [byte(240),159,140,182]
	':hotdog:': [byte(240),159,140,173]
	':hotel:': [byte(240),159,143,168]
	':hotsprings:': [byte(226),153,168]
	':hourglass:': [byte(226),140,155]
	':hourglass_flowing_sand:': [byte(226),143,179]
	':house:': [byte(240),159,143,160]
	':house_with_garden:': [byte(240),159,143,161]
	':houses:': [byte(240),159,143,152]
	':hugs:': [byte(240),159,164,151]
	':hungary:': [byte(240),159,135,173,240,159,135,186]
	':hushed:': [byte(240),159,152,175]
	':ice_cream:': [byte(240),159,141,168]
	':ice_cube:': [byte(240),159,167,138]
	':ice_hockey:': [byte(240),159,143,146]
	':ice_skate:': [byte(226),155,184]
	':icecream:': [byte(240),159,141,166]
	':iceland:': [byte(240),159,135,174,240,159,135,184]
	':id:': [byte(240),159,134,148]
	':ideograph_advantage:': [byte(240),159,137,144]
	':imp:': [byte(240),159,145,191]
	':inbox_tray:': [byte(240),159,147,165]
	':incoming_envelope:': [byte(240),159,147,168]
	':india:': [byte(240),159,135,174,240,159,135,179]
	':indonesia:': [byte(240),159,135,174,240,159,135,169]
	':infinity:': [byte(226),153,190]
	':information_desk_person:': [byte(240),159,146,129]
	':information_source:': [byte(226),132,185]
	':innocent:': [byte(240),159,152,135]
	':interrobang:': [byte(226),129,137]
	':iphone:': [byte(240),159,147,177]
	':iran:': [byte(240),159,135,174,240,159,135,183]
	':iraq:': [byte(240),159,135,174,240,159,135,182]
	':ireland:': [byte(240),159,135,174,240,159,135,170]
	':isle_of_man:': [byte(240),159,135,174,240,159,135,178]
	':israel:': [byte(240),159,135,174,240,159,135,177]
	':it:': [byte(240),159,135,174,240,159,135,185]
	':izakaya_lantern:': [byte(240),159,143,174]
	':jack_o_lantern:': [byte(240),159,142,131]
	':jamaica:': [byte(240),159,135,175,240,159,135,178]
	':japan:': [byte(240),159,151,190]
	':japanese_castle:': [byte(240),159,143,175]
	':japanese_goblin:': [byte(240),159,145,186]
	':japanese_ogre:': [byte(240),159,145,185]
	':jeans:': [byte(240),159,145,150]
	':jersey:': [byte(240),159,135,175,240,159,135,170]
	':jigsaw:': [byte(240),159,167,169]
	':jordan:': [byte(240),159,135,175,240,159,135,180]
	':joy:': [byte(240),159,152,130]
	':joy_cat:': [byte(240),159,152,185]
	':joystick:': [byte(240),159,149,185]
	':jp:': [byte(240),159,135,175,240,159,135,181]
	':judge:': [byte(240),159,167,145,226,154,150]
	':juggling_person:': [byte(240),159,164,185]
	':kaaba:': [byte(240),159,149,139]
	':kangaroo:': [byte(240),159,166,152]
	':kazakhstan:': [byte(240),159,135,176,240,159,135,191]
	':kenya:': [byte(240),159,135,176,240,159,135,170]
	':key:': [byte(240),159,148,145]
	':keyboard:': [byte(226),140,168]
	':keycap_ten:': [byte(240),159,148,159]
	':kick_scooter:': [byte(240),159,155,180]
	':kimono:': [byte(240),159,145,152]
	':kiribati:': [byte(240),159,135,176,240,159,135,174]
	':kiss:': [byte(240),159,146,139]
	':kissing:': [byte(240),159,152,151]
	':kissing_cat:': [byte(240),159,152,189]
	':kissing_closed_eyes:': [byte(240),159,152,154]
	':kissing_heart:': [byte(240),159,152,152]
	':kissing_smiling_eyes:': [byte(240),159,152,153]
	':kite:': [byte(240),159,170,129]
	':kiwi_fruit:': [byte(240),159,165,157]
	':kneeling_man:': [byte(240),159,167,142,226,153,130]
	':kneeling_person:': [byte(240),159,167,142]
	':kneeling_woman:': [byte(240),159,167,142,226,153,128]
	':knife:': [byte(240),159,148,170]
	':koala:': [byte(240),159,144,168]
	':koko:': [byte(240),159,136,129]
	':kosovo:': [byte(240),159,135,189,240,159,135,176]
	':kr:': [byte(240),159,135,176,240,159,135,183]
	':kuwait:': [byte(240),159,135,176,240,159,135,188]
	':kyrgyzstan:': [byte(240),159,135,176,240,159,135,172]
	':lab_coat:': [byte(240),159,165,188]
	':label:': [byte(240),159,143,183]
	':lacrosse:': [byte(240),159,165,141]
	':lantern:': [byte(240),159,143,174]
	':laos:': [byte(240),159,135,177,240,159,135,166]
	':large_blue_circle:': [byte(240),159,148,181]
	':large_blue_diamond:': [byte(240),159,148,183]
	':large_orange_diamond:': [byte(240),159,148,182]
	':last_quarter_moon:': [byte(240),159,140,151]
	':last_quarter_moon_with_face:': [byte(240),159,140,156]
	':latin_cross:': [byte(226),156,157]
	':latvia:': [byte(240),159,135,177,240,159,135,187]
	':laughing:': [byte(240),159,152,134]
	':leafy_green:': [byte(240),159,165,172]
	':leaves:': [byte(240),159,141,131]
	':lebanon:': [byte(240),159,135,177,240,159,135,167]
	':ledger:': [byte(240),159,147,146]
	':left_luggage:': [byte(240),159,155,133]
	':left_right_arrow:': [byte(226),134,148]
	':left_speech_bubble:': [byte(240),159,151,168]
	':leftwards_arrow_with_hook:': [byte(226),134,169]
	':leg:': [byte(240),159,166,181]
	':lemon:': [byte(240),159,141,139]
	':leo:': [byte(226),153,140]
	':leopard:': [byte(240),159,144,134]
	':lesotho:': [byte(240),159,135,177,240,159,135,184]
	':level_slider:': [byte(240),159,142,154]
	':liberia:': [byte(240),159,135,177,240,159,135,183]
	':libra:': [byte(226),153,142]
	':libya:': [byte(240),159,135,177,240,159,135,190]
	':liechtenstein:': [byte(240),159,135,177,240,159,135,174]
	':light_rail:': [byte(240),159,154,136]
	':link:': [byte(240),159,148,151]
	':lion:': [byte(240),159,166,129]
	':lips:': [byte(240),159,145,132]
	':lipstick:': [byte(240),159,146,132]
	':lithuania:': [byte(240),159,135,177,240,159,135,185]
	':lizard:': [byte(240),159,166,142]
	':llama:': [byte(240),159,166,153]
	':lobster:': [byte(240),159,166,158]
	':lock:': [byte(240),159,148,146]
	':lock_with_ink_pen:': [byte(240),159,148,143]
	':lollipop:': [byte(240),159,141,173]
	':loop:': [byte(226),158,191]
	':lotion_bottle:': [byte(240),159,167,180]
	':lotus_position:': [byte(240),159,167,152]
	':lotus_position_man:': [byte(240),159,167,152,226,153,130]
	':lotus_position_woman:': [byte(240),159,167,152,226,153,128]
	':loud_sound:': [byte(240),159,148,138]
	':loudspeaker:': [byte(240),159,147,162]
	':love_hotel:': [byte(240),159,143,169]
	':love_letter:': [byte(240),159,146,140]
	':love_you_gesture:': [byte(240),159,164,159]
	':low_brightness:': [byte(240),159,148,133]
	':luggage:': [byte(240),159,167,179]
	':luxembourg:': [byte(240),159,135,177,240,159,135,186]
	':lying_face:': [byte(240),159,164,165]
	':m:': [byte(226),147,130]
	':macau:': [byte(240),159,135,178,240,159,135,180]
	':macedonia:': [byte(240),159,135,178,240,159,135,176]
	':madagascar:': [byte(240),159,135,178,240,159,135,172]
	':mag:': [byte(240),159,148,141]
	':mag_right:': [byte(240),159,148,142]
	':mage:': [byte(240),159,167,153]
	':mage_man:': [byte(240),159,167,153,226,153,130]
	':mage_woman:': [byte(240),159,167,153,226,153,128]
	':magnet:': [byte(240),159,167,178]
	':mahjong:': [byte(240),159,128,132]
	':mailbox:': [byte(240),159,147,171]
	':mailbox_closed:': [byte(240),159,147,170]
	':mailbox_with_mail:': [byte(240),159,147,172]
	':mailbox_with_no_mail:': [byte(240),159,147,173]
	':malawi:': [byte(240),159,135,178,240,159,135,188]
	':malaysia:': [byte(240),159,135,178,240,159,135,190]
	':maldives:': [byte(240),159,135,178,240,159,135,187]
	':male_detective:': [byte(240),159,149,181,226,153,130]
	':male_sign:': [byte(226),153,130]
	':mali:': [byte(240),159,135,178,240,159,135,177]
	':malta:': [byte(240),159,135,178,240,159,135,185]
	':man:': [byte(240),159,145,168]
	':man_artist:': [byte(240),159,145,168,240,159,142,168]
	':man_astronaut:': [byte(240),159,145,168,240,159,154,128]
	':man_cartwheeling:': [byte(240),159,164,184,226,153,130]
	':man_cook:': [byte(240),159,145,168,240,159,141,179]
	':man_dancing:': [byte(240),159,149,186]
	':man_facepalming:': [byte(240),159,164,166,226,153,130]
	':man_factory_worker:': [byte(240),159,145,168,240,159,143,173]
	':man_farmer:': [byte(240),159,145,168,240,159,140,190]
	':man_firefighter:': [byte(240),159,145,168,240,159,154,146]
	':man_health_worker:': [byte(240),159,145,168,226,154,149]
	':man_in_manual_wheelchair:': [byte(240),159,145,168,240,159,166,189]
	':man_in_motorized_wheelchair:': [byte(240),159,145,168,240,159,166,188]
	':man_in_tuxedo:': [byte(240),159,164,181]
	':man_judge:': [byte(240),159,145,168,226,154,150]
	':man_juggling:': [byte(240),159,164,185,226,153,130]
	':man_mechanic:': [byte(240),159,145,168,240,159,148,167]
	':man_office_worker:': [byte(240),159,145,168,240,159,146,188]
	':man_pilot:': [byte(240),159,145,168,226,156,136]
	':man_playing_handball:': [byte(240),159,164,190,226,153,130]
	':man_playing_water_polo:': [byte(240),159,164,189,226,153,130]
	':man_scientist:': [byte(240),159,145,168,240,159,148,172]
	':man_shrugging:': [byte(240),159,164,183,226,153,130]
	':man_singer:': [byte(240),159,145,168,240,159,142,164]
	':man_student:': [byte(240),159,145,168,240,159,142,147]
	':man_teacher:': [byte(240),159,145,168,240,159,143,171]
	':man_technologist:': [byte(240),159,145,168,240,159,146,187]
	':man_with_gua_pi_mao:': [byte(240),159,145,178]
	':man_with_probing_cane:': [byte(240),159,145,168,240,159,166,175]
	':man_with_turban:': [byte(240),159,145,179,226,153,130]
	':mandarin:': [byte(240),159,141,138]
	':mango:': [byte(240),159,165,173]
	':mans_shoe:': [byte(240),159,145,158]
	':mantelpiece_clock:': [byte(240),159,149,176]
	':manual_wheelchair:': [byte(240),159,166,189]
	':maple_leaf:': [byte(240),159,141,129]
	':marshall_islands:': [byte(240),159,135,178,240,159,135,173]
	':martial_arts_uniform:': [byte(240),159,165,139]
	':martinique:': [byte(240),159,135,178,240,159,135,182]
	':mask:': [byte(240),159,152,183]
	':massage:': [byte(240),159,146,134]
	':massage_man:': [byte(240),159,146,134,226,153,130]
	':massage_woman:': [byte(240),159,146,134,226,153,128]
	':mate:': [byte(240),159,167,137]
	':mauritania:': [byte(240),159,135,178,240,159,135,183]
	':mauritius:': [byte(240),159,135,178,240,159,135,186]
	':mayotte:': [byte(240),159,135,190,240,159,135,185]
	':meat_on_bone:': [byte(240),159,141,150]
	':mechanic:': [byte(240),159,167,145,240,159,148,167]
	':mechanical_arm:': [byte(240),159,166,190]
	':mechanical_leg:': [byte(240),159,166,191]
	':medal_military:': [byte(240),159,142,150]
	':medal_sports:': [byte(240),159,143,133]
	':medical_symbol:': [byte(226),154,149]
	':mega:': [byte(240),159,147,163]
	':melon:': [byte(240),159,141,136]
	':memo:': [byte(240),159,147,157]
	':men_wrestling:': [byte(240),159,164,188,226,153,130]
	':menorah:': [byte(240),159,149,142]
	':mens:': [byte(240),159,154,185]
	':mermaid:': [byte(240),159,167,156,226,153,128]
	':merman:': [byte(240),159,167,156,226,153,130]
	':merperson:': [byte(240),159,167,156]
	':metal:': [byte(240),159,164,152]
	':metro:': [byte(240),159,154,135]
	':mexico:': [byte(240),159,135,178,240,159,135,189]
	':microbe:': [byte(240),159,166,160]
	':micronesia:': [byte(240),159,135,171,240,159,135,178]
	':microphone:': [byte(240),159,142,164]
	':microscope:': [byte(240),159,148,172]
	':middle_finger:': [byte(240),159,150,149]
	':milk_glass:': [byte(240),159,165,155]
	':milky_way:': [byte(240),159,140,140]
	':minibus:': [byte(240),159,154,144]
	':minidisc:': [byte(240),159,146,189]
	':mobile_phone_off:': [byte(240),159,147,180]
	':moldova:': [byte(240),159,135,178,240,159,135,169]
	':monaco:': [byte(240),159,135,178,240,159,135,168]
	':money_mouth_face:': [byte(240),159,164,145]
	':money_with_wings:': [byte(240),159,146,184]
	':moneybag:': [byte(240),159,146,176]
	':mongolia:': [byte(240),159,135,178,240,159,135,179]
	':monkey:': [byte(240),159,144,146]
	':monkey_face:': [byte(240),159,144,181]
	':monocle_face:': [byte(240),159,167,144]
	':monorail:': [byte(240),159,154,157]
	':montenegro:': [byte(240),159,135,178,240,159,135,170]
	':montserrat:': [byte(240),159,135,178,240,159,135,184]
	':moon:': [byte(240),159,140,148]
	':moon_cake:': [byte(240),159,165,174]
	':morocco:': [byte(240),159,135,178,240,159,135,166]
	':mortar_board:': [byte(240),159,142,147]
	':mosque:': [byte(240),159,149,140]
	':mosquito:': [byte(240),159,166,159]
	':motor_boat:': [byte(240),159,155,165]
	':motor_scooter:': [byte(240),159,155,181]
	':motorcycle:': [byte(240),159,143,141]
	':motorized_wheelchair:': [byte(240),159,166,188]
	':motorway:': [byte(240),159,155,163]
	':mount_fuji:': [byte(240),159,151,187]
	':mountain:': [byte(226),155,176]
	':mountain_bicyclist:': [byte(240),159,154,181]
	':mountain_biking_man:': [byte(240),159,154,181,226,153,130]
	':mountain_biking_woman:': [byte(240),159,154,181,226,153,128]
	':mountain_cableway:': [byte(240),159,154,160]
	':mountain_railway:': [byte(240),159,154,158]
	':mountain_snow:': [byte(240),159,143,148]
	':mouse:': [byte(240),159,144,173]
	':mouse2:': [byte(240),159,144,129]
	':movie_camera:': [byte(240),159,142,165]
	':moyai:': [byte(240),159,151,191]
	':mozambique:': [byte(240),159,135,178,240,159,135,191]
	':mrs_claus:': [byte(240),159,164,182]
	':muscle:': [byte(240),159,146,170]
	':mushroom:': [byte(240),159,141,132]
	':musical_keyboard:': [byte(240),159,142,185]
	':musical_note:': [byte(240),159,142,181]
	':musical_score:': [byte(240),159,142,188]
	':mute:': [byte(240),159,148,135]
	':myanmar:': [byte(240),159,135,178,240,159,135,178]
	':nail_care:': [byte(240),159,146,133]
	':name_badge:': [byte(240),159,147,155]
	':namibia:': [byte(240),159,135,179,240,159,135,166]
	':national_park:': [byte(240),159,143,158]
	':nauru:': [byte(240),159,135,179,240,159,135,183]
	':nauseated_face:': [byte(240),159,164,162]
	':nazar_amulet:': [byte(240),159,167,191]
	':necktie:': [byte(240),159,145,148]
	':negative_squared_cross_mark:': [byte(226),157,142]
	':nepal:': [byte(240),159,135,179,240,159,135,181]
	':nerd_face:': [byte(240),159,164,147]
	':netherlands:': [byte(240),159,135,179,240,159,135,177]
	':neutral_face:': [byte(240),159,152,144]
	':new:': [byte(240),159,134,149]
	':new_caledonia:': [byte(240),159,135,179,240,159,135,168]
	':new_moon:': [byte(240),159,140,145]
	':new_moon_with_face:': [byte(240),159,140,154]
	':new_zealand:': [byte(240),159,135,179,240,159,135,191]
	':newspaper:': [byte(240),159,147,176]
	':newspaper_roll:': [byte(240),159,151,158]
	':next_track_button:': [byte(226),143,173]
	':ng:': [byte(240),159,134,150]
	':ng_man:': [byte(240),159,153,133,226,153,130]
	':ng_woman:': [byte(240),159,153,133,226,153,128]
	':nicaragua:': [byte(240),159,135,179,240,159,135,174]
	':niger:': [byte(240),159,135,179,240,159,135,170]
	':nigeria:': [byte(240),159,135,179,240,159,135,172]
	':night_with_stars:': [byte(240),159,140,131]
	':nine:': [byte(57),226,131,163]
	':niue:': [byte(240),159,135,179,240,159,135,186]
	':no_bell:': [byte(240),159,148,149]
	':no_bicycles:': [byte(240),159,154,179]
	':no_entry:': [byte(226),155,148]
	':no_entry_sign:': [byte(240),159,154,171]
	':no_good:': [byte(240),159,153,133]
	':no_good_man:': [byte(240),159,153,133,226,153,130]
	':no_good_woman:': [byte(240),159,153,133,226,153,128]
	':no_mobile_phones:': [byte(240),159,147,181]
	':no_mouth:': [byte(240),159,152,182]
	':no_pedestrians:': [byte(240),159,154,183]
	':no_smoking:': [byte(240),159,154,173]
	':non-potable_water:': [byte(240),159,154,177]
	':norfolk_island:': [byte(240),159,135,179,240,159,135,171]
	':north_korea:': [byte(240),159,135,176,240,159,135,181]
	':northern_mariana_islands:': [byte(240),159,135,178,240,159,135,181]
	':norway:': [byte(240),159,135,179,240,159,135,180]
	':nose:': [byte(240),159,145,131]
	':notebook:': [byte(240),159,147,147]
	':notebook_with_decorative_cover:': [byte(240),159,147,148]
	':notes:': [byte(240),159,142,182]
	':nut_and_bolt:': [byte(240),159,148,169]
	':o:': [byte(226),173,149]
	':o2:': [byte(240),159,133,190]
	':ocean:': [byte(240),159,140,138]
	':octopus:': [byte(240),159,144,153]
	':oden:': [byte(240),159,141,162]
	':office:': [byte(240),159,143,162]
	':office_worker:': [byte(240),159,167,145,240,159,146,188]
	':oil_drum:': [byte(240),159,155,162]
	':ok:': [byte(240),159,134,151]
	':ok_hand:': [byte(240),159,145,140]
	':ok_man:': [byte(240),159,153,134,226,153,130]
	':ok_person:': [byte(240),159,153,134]
	':ok_woman:': [byte(240),159,153,134,226,153,128]
	':old_key:': [byte(240),159,151,157]
	':older_adult:': [byte(240),159,167,147]
	':older_man:': [byte(240),159,145,180]
	':older_woman:': [byte(240),159,145,181]
	':om:': [byte(240),159,149,137]
	':oman:': [byte(240),159,135,180,240,159,135,178]
	':on:': [byte(240),159,148,155]
	':oncoming_automobile:': [byte(240),159,154,152]
	':oncoming_bus:': [byte(240),159,154,141]
	':oncoming_police_car:': [byte(240),159,154,148]
	':oncoming_taxi:': [byte(240),159,154,150]
	':one:': [byte(49),226,131,163]
	':one_piece_swimsuit:': [byte(240),159,169,177]
	':onion:': [byte(240),159,167,133]
	':open_book:': [byte(240),159,147,150]
	':open_file_folder:': [byte(240),159,147,130]
	':open_hands:': [byte(240),159,145,144]
	':open_mouth:': [byte(240),159,152,174]
	':open_umbrella:': [byte(226),152,130]
	':ophiuchus:': [byte(226),155,142]
	':orange:': [byte(240),159,141,138]
	':orange_book:': [byte(240),159,147,153]
	':orange_circle:': [byte(240),159,159,160]
	':orange_heart:': [byte(240),159,167,161]
	':orange_square:': [byte(240),159,159,167]
	':orangutan:': [byte(240),159,166,167]
	':orthodox_cross:': [byte(226),152,166]
	':otter:': [byte(240),159,166,166]
	':outbox_tray:': [byte(240),159,147,164]
	':owl:': [byte(240),159,166,137]
	':ox:': [byte(240),159,144,130]
	':oyster:': [byte(240),159,166,170]
	':package:': [byte(240),159,147,166]
	':page_facing_up:': [byte(240),159,147,132]
	':page_with_curl:': [byte(240),159,147,131]
	':pager:': [byte(240),159,147,159]
	':paintbrush:': [byte(240),159,150,140]
	':pakistan:': [byte(240),159,135,181,240,159,135,176]
	':palau:': [byte(240),159,135,181,240,159,135,188]
	':palestinian_territories:': [byte(240),159,135,181,240,159,135,184]
	':palm_tree:': [byte(240),159,140,180]
	':palms_up_together:': [byte(240),159,164,178]
	':panama:': [byte(240),159,135,181,240,159,135,166]
	':pancakes:': [byte(240),159,165,158]
	':panda_face:': [byte(240),159,144,188]
	':paperclip:': [byte(240),159,147,142]
	':paperclips:': [byte(240),159,150,135]
	':papua_new_guinea:': [byte(240),159,135,181,240,159,135,172]
	':parachute:': [byte(240),159,170,130]
	':paraguay:': [byte(240),159,135,181,240,159,135,190]
	':parasol_on_ground:': [byte(226),155,177]
	':parking:': [byte(240),159,133,191]
	':parrot:': [byte(240),159,166,156]
	':part_alternation_mark:': [byte(227),128,189]
	':partly_sunny:': [byte(226),155,133]
	':partying_face:': [byte(240),159,165,179]
	':passenger_ship:': [byte(240),159,155,179]
	':passport_control:': [byte(240),159,155,130]
	':pause_button:': [byte(226),143,184]
	':paw_prints:': [byte(240),159,144,190]
	':peace_symbol:': [byte(226),152,174]
	':peach:': [byte(240),159,141,145]
	':peacock:': [byte(240),159,166,154]
	':peanuts:': [byte(240),159,165,156]
	':pear:': [byte(240),159,141,144]
	':pen:': [byte(240),159,150,138]
	':pencil:': [byte(240),159,147,157]
	':pencil2:': [byte(226),156,143]
	':penguin:': [byte(240),159,144,167]
	':pensive:': [byte(240),159,152,148]
	':people_holding_hands:': [byte(240),159,167,145,240,159,164,157,240,159,167,145]
	':performing_arts:': [byte(240),159,142,173]
	':persevere:': [byte(240),159,152,163]
	':person_bald:': [byte(240),159,167,145,240,159,166,178]
	':person_curly_hair:': [byte(240),159,167,145,240,159,166,177]
	':person_fencing:': [byte(240),159,164,186]
	':person_in_manual_wheelchair:': [byte(240),159,167,145,240,159,166,189]
	':person_in_motorized_wheelchair:': [byte(240),159,167,145,240,159,166,188]
	':person_red_hair:': [byte(240),159,167,145,240,159,166,176]
	':person_white_hair:': [byte(240),159,167,145,240,159,166,179]
	':person_with_probing_cane:': [byte(240),159,167,145,240,159,166,175]
	':person_with_turban:': [byte(240),159,145,179]
	':peru:': [byte(240),159,135,181,240,159,135,170]
	':petri_dish:': [byte(240),159,167,171]
	':philippines:': [byte(240),159,135,181,240,159,135,173]
	':phone:': [byte(226),152,142]
	':pick:': [byte(226),155,143]
	':pie:': [byte(240),159,165,167]
	':pig:': [byte(240),159,144,183]
	':pig2:': [byte(240),159,144,150]
	':pig_nose:': [byte(240),159,144,189]
	':pill:': [byte(240),159,146,138]
	':pilot:': [byte(240),159,167,145,226,156,136]
	':pinching_hand:': [byte(240),159,164,143]
	':pineapple:': [byte(240),159,141,141]
	':ping_pong:': [byte(240),159,143,147]
	':pirate_flag:': [byte(240),159,143,180,226,152,160]
	':pisces:': [byte(226),153,147]
	':pitcairn_islands:': [byte(240),159,135,181,240,159,135,179]
	':pizza:': [byte(240),159,141,149]
	':place_of_worship:': [byte(240),159,155,144]
	':plate_with_cutlery:': [byte(240),159,141,189]
	':play_or_pause_button:': [byte(226),143,175]
	':pleading_face:': [byte(240),159,165,186]
	':point_down:': [byte(240),159,145,135]
	':point_left:': [byte(240),159,145,136]
	':point_right:': [byte(240),159,145,137]
	':point_up:': [byte(226),152,157]
	':point_up_2:': [byte(240),159,145,134]
	':poland:': [byte(240),159,135,181,240,159,135,177]
	':police_car:': [byte(240),159,154,147]
	':police_officer:': [byte(240),159,145,174]
	':policeman:': [byte(240),159,145,174,226,153,130]
	':policewoman:': [byte(240),159,145,174,226,153,128]
	':poodle:': [byte(240),159,144,169]
	':poop:': [byte(240),159,146,169]
	':popcorn:': [byte(240),159,141,191]
	':portugal:': [byte(240),159,135,181,240,159,135,185]
	':post_office:': [byte(240),159,143,163]
	':postal_horn:': [byte(240),159,147,175]
	':postbox:': [byte(240),159,147,174]
	':potable_water:': [byte(240),159,154,176]
	':potato:': [byte(240),159,165,148]
	':pouch:': [byte(240),159,145,157]
	':poultry_leg:': [byte(240),159,141,151]
	':pound:': [byte(240),159,146,183]
	':pout:': [byte(240),159,152,161]
	':pouting_cat:': [byte(240),159,152,190]
	':pouting_face:': [byte(240),159,153,142]
	':pouting_man:': [byte(240),159,153,142,226,153,130]
	':pouting_woman:': [byte(240),159,153,142,226,153,128]
	':pray:': [byte(240),159,153,143]
	':prayer_beads:': [byte(240),159,147,191]
	':pregnant_woman:': [byte(240),159,164,176]
	':pretzel:': [byte(240),159,165,168]
	':previous_track_button:': [byte(226),143,174]
	':prince:': [byte(240),159,164,180]
	':princess:': [byte(240),159,145,184]
	':printer:': [byte(240),159,150,168]
	':probing_cane:': [byte(240),159,166,175]
	':puerto_rico:': [byte(240),159,135,181,240,159,135,183]
	':punch:': [byte(240),159,145,138]
	':purple_circle:': [byte(240),159,159,163]
	':purple_heart:': [byte(240),159,146,156]
	':purple_square:': [byte(240),159,159,170]
	':purse:': [byte(240),159,145,155]
	':pushpin:': [byte(240),159,147,140]
	':put_litter_in_its_place:': [byte(240),159,154,174]
	':qatar:': [byte(240),159,135,182,240,159,135,166]
	':question:': [byte(226),157,147]
	':rabbit:': [byte(240),159,144,176]
	':rabbit2:': [byte(240),159,144,135]
	':raccoon:': [byte(240),159,166,157]
	':racehorse:': [byte(240),159,144,142]
	':racing_car:': [byte(240),159,143,142]
	':radio:': [byte(240),159,147,187]
	':radio_button:': [byte(240),159,148,152]
	':radioactive:': [byte(226),152,162]
	':rage:': [byte(240),159,152,161]
	':railway_car:': [byte(240),159,154,131]
	':railway_track:': [byte(240),159,155,164]
	':rainbow:': [byte(240),159,140,136]
	':rainbow_flag:': [byte(240),159,143,179,240,159,140,136]
	':raised_back_of_hand:': [byte(240),159,164,154]
	':raised_eyebrow:': [byte(240),159,164,168]
	':raised_hand:': [byte(226),156,139]
	':raised_hand_with_fingers_splayed:': [byte(240),159,150,144]
	':raised_hands:': [byte(240),159,153,140]
	':raising_hand:': [byte(240),159,153,139]
	':raising_hand_man:': [byte(240),159,153,139,226,153,130]
	':raising_hand_woman:': [byte(240),159,153,139,226,153,128]
	':ram:': [byte(240),159,144,143]
	':ramen:': [byte(240),159,141,156]
	':rat:': [byte(240),159,144,128]
	':razor:': [byte(240),159,170,146]
	':receipt:': [byte(240),159,167,190]
	':record_button:': [byte(226),143,186]
	':recycle:': [byte(226),153,187]
	':red_car:': [byte(240),159,154,151]
	':red_circle:': [byte(240),159,148,180]
	':red_envelope:': [byte(240),159,167,167]
	':red_haired_man:': [byte(240),159,145,168,240,159,166,176]
	':red_haired_woman:': [byte(240),159,145,169,240,159,166,176]
	':red_square:': [byte(240),159,159,165]
	':registered:': [byte(194),174]
	':relaxed:': [byte(226),152,186]
	':relieved:': [byte(240),159,152,140]
	':reminder_ribbon:': [byte(240),159,142,151]
	':repeat:': [byte(240),159,148,129]
	':repeat_one:': [byte(240),159,148,130]
	':rescue_worker_helmet:': [byte(226),155,145]
	':restroom:': [byte(240),159,154,187]
	':reunion:': [byte(240),159,135,183,240,159,135,170]
	':revolving_hearts:': [byte(240),159,146,158]
	':rewind:': [byte(226),143,170]
	':rhinoceros:': [byte(240),159,166,143]
	':ribbon:': [byte(240),159,142,128]
	':rice:': [byte(240),159,141,154]
	':rice_ball:': [byte(240),159,141,153]
	':rice_cracker:': [byte(240),159,141,152]
	':rice_scene:': [byte(240),159,142,145]
	':right_anger_bubble:': [byte(240),159,151,175]
	':ring:': [byte(240),159,146,141]
	':ringed_planet:': [byte(240),159,170,144]
	':robot:': [byte(240),159,164,150]
	':rocket:': [byte(240),159,154,128]
	':rofl:': [byte(240),159,164,163]
	':roll_eyes:': [byte(240),159,153,132]
	':roll_of_paper:': [byte(240),159,167,187]
	':roller_coaster:': [byte(240),159,142,162]
	':romania:': [byte(240),159,135,183,240,159,135,180]
	':rooster:': [byte(240),159,144,147]
	':rose:': [byte(240),159,140,185]
	':rosette:': [byte(240),159,143,181]
	':rotating_light:': [byte(240),159,154,168]
	':round_pushpin:': [byte(240),159,147,141]
	':rowboat:': [byte(240),159,154,163]
	':rowing_man:': [byte(240),159,154,163,226,153,130]
	':rowing_woman:': [byte(240),159,154,163,226,153,128]
	':ru:': [byte(240),159,135,183,240,159,135,186]
	':rugby_football:': [byte(240),159,143,137]
	':runner:': [byte(240),159,143,131]
	':running:': [byte(240),159,143,131]
	':running_man:': [byte(240),159,143,131,226,153,130]
	':running_shirt_with_sash:': [byte(240),159,142,189]
	':running_woman:': [byte(240),159,143,131,226,153,128]
	':rwanda:': [byte(240),159,135,183,240,159,135,188]
	':sa:': [byte(240),159,136,130]
	':safety_pin:': [byte(240),159,167,183]
	':safety_vest:': [byte(240),159,166,186]
	':sagittarius:': [byte(226),153,144]
	':sailboat:': [byte(226),155,181]
	':sake:': [byte(240),159,141,182]
	':salt:': [byte(240),159,167,130]
	':samoa:': [byte(240),159,135,188,240,159,135,184]
	':san_marino:': [byte(240),159,135,184,240,159,135,178]
	':sandal:': [byte(240),159,145,161]
	':sandwich:': [byte(240),159,165,170]
	':santa:': [byte(240),159,142,133]
	':sao_tome_principe:': [byte(240),159,135,184,240,159,135,185]
	':sari:': [byte(240),159,165,187]
	':sassy_man:': [byte(240),159,146,129,226,153,130]
	':sassy_woman:': [byte(240),159,146,129,226,153,128]
	':satellite:': [byte(240),159,147,161]
	':satisfied:': [byte(240),159,152,134]
	':saudi_arabia:': [byte(240),159,135,184,240,159,135,166]
	':sauna_man:': [byte(240),159,167,150,226,153,130]
	':sauna_person:': [byte(240),159,167,150]
	':sauna_woman:': [byte(240),159,167,150,226,153,128]
	':sauropod:': [byte(240),159,166,149]
	':saxophone:': [byte(240),159,142,183]
	':scarf:': [byte(240),159,167,163]
	':school:': [byte(240),159,143,171]
	':school_satchel:': [byte(240),159,142,146]
	':scientist:': [byte(240),159,167,145,240,159,148,172]
	':scissors:': [byte(226),156,130]
	':scorpion:': [byte(240),159,166,130]
	':scorpius:': [byte(226),153,143]
	':scotland:': [byte(240),159,143,180,243,160,129,167,243,160,129,162,243,160,129,179,243,160,129,163,243,160,129,180,243,160,129,191]
	':scream:': [byte(240),159,152,177]
	':scream_cat:': [byte(240),159,153,128]
	':scroll:': [byte(240),159,147,156]
	':seat:': [byte(240),159,146,186]
	':secret:': [byte(227),138,153]
	':see_no_evil:': [byte(240),159,153,136]
	':seedling:': [byte(240),159,140,177]
	':selfie:': [byte(240),159,164,179]
	':senegal:': [byte(240),159,135,184,240,159,135,179]
	':serbia:': [byte(240),159,135,183,240,159,135,184]
	':service_dog:': [byte(240),159,144,149,240,159,166,186]
	':seven:': [byte(55),226,131,163]
	':seychelles:': [byte(240),159,135,184,240,159,135,168]
	':shallow_pan_of_food:': [byte(240),159,165,152]
	':shamrock:': [byte(226),152,152]
	':shark:': [byte(240),159,166,136]
	':shaved_ice:': [byte(240),159,141,167]
	':sheep:': [byte(240),159,144,145]
	':shell:': [byte(240),159,144,154]
	':shield:': [byte(240),159,155,161]
	':shinto_shrine:': [byte(226),155,169]
	':ship:': [byte(240),159,154,162]
	':shirt:': [byte(240),159,145,149]
	':shit:': [byte(240),159,146,169]
	':shoe:': [byte(240),159,145,158]
	':shopping:': [byte(240),159,155,141]
	':shopping_cart:': [byte(240),159,155,146]
	':shorts:': [byte(240),159,169,179]
	':shower:': [byte(240),159,154,191]
	':shrimp:': [byte(240),159,166,144]
	':shrug:': [byte(240),159,164,183]
	':shushing_face:': [byte(240),159,164,171]
	':sierra_leone:': [byte(240),159,135,184,240,159,135,177]
	':signal_strength:': [byte(240),159,147,182]
	':singapore:': [byte(240),159,135,184,240,159,135,172]
	':singer:': [byte(240),159,167,145,240,159,142,164]
	':sint_maarten:': [byte(240),159,135,184,240,159,135,189]
	':six:': [byte(54),226,131,163]
	':six_pointed_star:': [byte(240),159,148,175]
	':skateboard:': [byte(240),159,155,185]
	':ski:': [byte(240),159,142,191]
	':skier:': [byte(226),155,183]
	':skull:': [byte(240),159,146,128]
	':skull_and_crossbones:': [byte(226),152,160]
	':skunk:': [byte(240),159,166,168]
	':sled:': [byte(240),159,155,183]
	':sleeping:': [byte(240),159,152,180]
	':sleeping_bed:': [byte(240),159,155,140]
	':sleepy:': [byte(240),159,152,170]
	':slightly_frowning_face:': [byte(240),159,153,129]
	':slightly_smiling_face:': [byte(240),159,153,130]
	':slot_machine:': [byte(240),159,142,176]
	':sloth:': [byte(240),159,166,165]
	':slovakia:': [byte(240),159,135,184,240,159,135,176]
	':slovenia:': [byte(240),159,135,184,240,159,135,174]
	':small_airplane:': [byte(240),159,155,169]
	':small_blue_diamond:': [byte(240),159,148,185]
	':small_orange_diamond:': [byte(240),159,148,184]
	':small_red_triangle:': [byte(240),159,148,186]
	':small_red_triangle_down:': [byte(240),159,148,187]
	':smile:': [byte(240),159,152,132]
	':smile_cat:': [byte(240),159,152,184]
	':smiley:': [byte(240),159,152,131]
	':smiley_cat:': [byte(240),159,152,186]
	':smiling_face_with_three_hearts:': [byte(240),159,165,176]
	':smiling_imp:': [byte(240),159,152,136]
	':smirk:': [byte(240),159,152,143]
	':smirk_cat:': [byte(240),159,152,188]
	':smoking:': [byte(240),159,154,172]
	':snail:': [byte(240),159,144,140]
	':snake:': [byte(240),159,144,141]
	':sneezing_face:': [byte(240),159,164,167]
	':snowboarder:': [byte(240),159,143,130]
	':snowflake:': [byte(226),157,132]
	':snowman:': [byte(226),155,132]
	':snowman_with_snow:': [byte(226),152,131]
	':soap:': [byte(240),159,167,188]
	':sob:': [byte(240),159,152,173]
	':soccer:': [byte(226),154,189]
	':socks:': [byte(240),159,167,166]
	':softball:': [byte(240),159,165,142]
	':solomon_islands:': [byte(240),159,135,184,240,159,135,167]
	':somalia:': [byte(240),159,135,184,240,159,135,180]
	':soon:': [byte(240),159,148,156]
	':sos:': [byte(240),159,134,152]
	':sound:': [byte(240),159,148,137]
	':south_africa:': [byte(240),159,135,191,240,159,135,166]
	':south_georgia_south_sandwich_islands:': [byte(240),159,135,172,240,159,135,184]
	':south_sudan:': [byte(240),159,135,184,240,159,135,184]
	':space_invader:': [byte(240),159,145,190]
	':spades:': [byte(226),153,160]
	':spaghetti:': [byte(240),159,141,157]
	':sparkle:': [byte(226),157,135]
	':sparkler:': [byte(240),159,142,135]
	':sparkles:': [byte(226),156,168]
	':sparkling_heart:': [byte(240),159,146,150]
	':speak_no_evil:': [byte(240),159,153,138]
	':speaker:': [byte(240),159,148,136]
	':speaking_head:': [byte(240),159,151,163]
	':speech_balloon:': [byte(240),159,146,172]
	':speedboat:': [byte(240),159,154,164]
	':spider:': [byte(240),159,149,183]
	':spider_web:': [byte(240),159,149,184]
	':spiral_calendar:': [byte(240),159,151,147]
	':spiral_notepad:': [byte(240),159,151,146]
	':sponge:': [byte(240),159,167,189]
	':spoon:': [byte(240),159,165,132]
	':squid:': [byte(240),159,166,145]
	':sri_lanka:': [byte(240),159,135,177,240,159,135,176]
	':st_barthelemy:': [byte(240),159,135,167,240,159,135,177]
	':st_helena:': [byte(240),159,135,184,240,159,135,173]
	':st_kitts_nevis:': [byte(240),159,135,176,240,159,135,179]
	':st_lucia:': [byte(240),159,135,177,240,159,135,168]
	':st_martin:': [byte(240),159,135,178,240,159,135,171]
	':st_pierre_miquelon:': [byte(240),159,135,181,240,159,135,178]
	':st_vincent_grenadines:': [byte(240),159,135,187,240,159,135,168]
	':stadium:': [byte(240),159,143,159]
	':standing_man:': [byte(240),159,167,141,226,153,130]
	':standing_person:': [byte(240),159,167,141]
	':standing_woman:': [byte(240),159,167,141,226,153,128]
	':star:': [byte(226),173,144]
	':star2:': [byte(240),159,140,159]
	':star_and_crescent:': [byte(226),152,170]
	':star_of_david:': [byte(226),156,161]
	':star_struck:': [byte(240),159,164,169]
	':stars:': [byte(240),159,140,160]
	':station:': [byte(240),159,154,137]
	':statue_of_liberty:': [byte(240),159,151,189]
	':steam_locomotive:': [byte(240),159,154,130]
	':stethoscope:': [byte(240),159,169,186]
	':stew:': [byte(240),159,141,178]
	':stop_button:': [byte(226),143,185]
	':stop_sign:': [byte(240),159,155,145]
	':stopwatch:': [byte(226),143,177]
	':straight_ruler:': [byte(240),159,147,143]
	':strawberry:': [byte(240),159,141,147]
	':stuck_out_tongue:': [byte(240),159,152,155]
	':stuck_out_tongue_closed_eyes:': [byte(240),159,152,157]
	':stuck_out_tongue_winking_eye:': [byte(240),159,152,156]
	':student:': [byte(240),159,167,145,240,159,142,147]
	':studio_microphone:': [byte(240),159,142,153]
	':stuffed_flatbread:': [byte(240),159,165,153]
	':sudan:': [byte(240),159,135,184,240,159,135,169]
	':sun_behind_large_cloud:': [byte(240),159,140,165]
	':sun_behind_rain_cloud:': [byte(240),159,140,166]
	':sun_behind_small_cloud:': [byte(240),159,140,164]
	':sun_with_face:': [byte(240),159,140,158]
	':sunflower:': [byte(240),159,140,187]
	':sunglasses:': [byte(240),159,152,142]
	':sunny:': [byte(226),152,128]
	':sunrise:': [byte(240),159,140,133]
	':sunrise_over_mountains:': [byte(240),159,140,132]
	':superhero:': [byte(240),159,166,184]
	':superhero_man:': [byte(240),159,166,184,226,153,130]
	':superhero_woman:': [byte(240),159,166,184,226,153,128]
	':supervillain:': [byte(240),159,166,185]
	':supervillain_man:': [byte(240),159,166,185,226,153,130]
	':supervillain_woman:': [byte(240),159,166,185,226,153,128]
	':surfer:': [byte(240),159,143,132]
	':surfing_man:': [byte(240),159,143,132,226,153,130]
	':surfing_woman:': [byte(240),159,143,132,226,153,128]
	':suriname:': [byte(240),159,135,184,240,159,135,183]
	':sushi:': [byte(240),159,141,163]
	':suspension_railway:': [byte(240),159,154,159]
	':svalbard_jan_mayen:': [byte(240),159,135,184,240,159,135,175]
	':swan:': [byte(240),159,166,162]
	':swaziland:': [byte(240),159,135,184,240,159,135,191]
	':sweat:': [byte(240),159,152,147]
	':sweat_drops:': [byte(240),159,146,166]
	':sweat_smile:': [byte(240),159,152,133]
	':sweden:': [byte(240),159,135,184,240,159,135,170]
	':sweet_potato:': [byte(240),159,141,160]
	':swim_brief:': [byte(240),159,169,178]
	':swimmer:': [byte(240),159,143,138]
	':swimming_man:': [byte(240),159,143,138,226,153,130]
	':swimming_woman:': [byte(240),159,143,138,226,153,128]
	':switzerland:': [byte(240),159,135,168,240,159,135,173]
	':symbols:': [byte(240),159,148,163]
	':synagogue:': [byte(240),159,149,141]
	':syria:': [byte(240),159,135,184,240,159,135,190]
	':syringe:': [byte(240),159,146,137]
	':t-rex:': [byte(240),159,166,150]
	':taco:': [byte(240),159,140,174]
	':tada:': [byte(240),159,142,137]
	':taiwan:': [byte(240),159,135,185,240,159,135,188]
	':tajikistan:': [byte(240),159,135,185,240,159,135,175]
	':takeout_box:': [byte(240),159,165,161]
	':tanabata_tree:': [byte(240),159,142,139]
	':tangerine:': [byte(240),159,141,138]
	':tanzania:': [byte(240),159,135,185,240,159,135,191]
	':taurus:': [byte(226),153,137]
	':taxi:': [byte(240),159,154,149]
	':tea:': [byte(240),159,141,181]
	':teacher:': [byte(240),159,167,145,240,159,143,171]
	':technologist:': [byte(240),159,167,145,240,159,146,187]
	':teddy_bear:': [byte(240),159,167,184]
	':telephone:': [byte(226),152,142]
	':telephone_receiver:': [byte(240),159,147,158]
	':telescope:': [byte(240),159,148,173]
	':tennis:': [byte(240),159,142,190]
	':tent:': [byte(226),155,186]
	':test_tube:': [byte(240),159,167,170]
	':thailand:': [byte(240),159,135,185,240,159,135,173]
	':thermometer:': [byte(240),159,140,161]
	':thinking:': [byte(240),159,164,148]
	':thought_balloon:': [byte(240),159,146,173]
	':thread:': [byte(240),159,167,181]
	':three:': [byte(51),226,131,163]
	':thumbsdown:': [byte(240),159,145,142]
	':thumbsup:': [byte(240),159,145,141]
	':ticket:': [byte(240),159,142,171]
	':tickets:': [byte(240),159,142,159]
	':tiger:': [byte(240),159,144,175]
	':tiger2:': [byte(240),159,144,133]
	':timer_clock:': [byte(226),143,178]
	':timor_leste:': [byte(240),159,135,185,240,159,135,177]
	':tipping_hand_man:': [byte(240),159,146,129,226,153,130]
	':tipping_hand_person:': [byte(240),159,146,129]
	':tipping_hand_woman:': [byte(240),159,146,129,226,153,128]
	':tired_face:': [byte(240),159,152,171]
	':tm:': [byte(226),132,162]
	':togo:': [byte(240),159,135,185,240,159,135,172]
	':toilet:': [byte(240),159,154,189]
	':tokelau:': [byte(240),159,135,185,240,159,135,176]
	':tokyo_tower:': [byte(240),159,151,188]
	':tomato:': [byte(240),159,141,133]
	':tonga:': [byte(240),159,135,185,240,159,135,180]
	':tongue:': [byte(240),159,145,133]
	':toolbox:': [byte(240),159,167,176]
	':tooth:': [byte(240),159,166,183]
	':top:': [byte(240),159,148,157]
	':tophat:': [byte(240),159,142,169]
	':tornado:': [byte(240),159,140,170]
	':tr:': [byte(240),159,135,185,240,159,135,183]
	':trackball:': [byte(240),159,150,178]
	':tractor:': [byte(240),159,154,156]
	':traffic_light:': [byte(240),159,154,165]
	':train:': [byte(240),159,154,139]
	':train2:': [byte(240),159,154,134]
	':tram:': [byte(240),159,154,138]
	':triangular_flag_on_post:': [byte(240),159,154,169]
	':triangular_ruler:': [byte(240),159,147,144]
	':trident:': [byte(240),159,148,177]
	':trinidad_tobago:': [byte(240),159,135,185,240,159,135,185]
	':tristan_da_cunha:': [byte(240),159,135,185,240,159,135,166]
	':triumph:': [byte(240),159,152,164]
	':trolleybus:': [byte(240),159,154,142]
	':trophy:': [byte(240),159,143,134]
	':tropical_drink:': [byte(240),159,141,185]
	':tropical_fish:': [byte(240),159,144,160]
	':truck:': [byte(240),159,154,154]
	':trumpet:': [byte(240),159,142,186]
	':tshirt:': [byte(240),159,145,149]
	':tulip:': [byte(240),159,140,183]
	':tumbler_glass:': [byte(240),159,165,131]
	':tunisia:': [byte(240),159,135,185,240,159,135,179]
	':turkey:': [byte(240),159,166,131]
	':turkmenistan:': [byte(240),159,135,185,240,159,135,178]
	':turks_caicos_islands:': [byte(240),159,135,185,240,159,135,168]
	':turtle:': [byte(240),159,144,162]
	':tuvalu:': [byte(240),159,135,185,240,159,135,187]
	':tv:': [byte(240),159,147,186]
	':twisted_rightwards_arrows:': [byte(240),159,148,128]
	':two:': [byte(50),226,131,163]
	':two_hearts:': [byte(240),159,146,149]
	':two_men_holding_hands:': [byte(240),159,145,172]
	':two_women_holding_hands:': [byte(240),159,145,173]
	':u5272:': [byte(240),159,136,185]
	':u5408:': [byte(240),159,136,180]
	':u55b6:': [byte(240),159,136,186]
	':u6307:': [byte(240),159,136,175]
	':u6708:': [byte(240),159,136,183]
	':u6709:': [byte(240),159,136,182]
	':u6e80:': [byte(240),159,136,181]
	':u7121:': [byte(240),159,136,154]
	':u7533:': [byte(240),159,136,184]
	':u7981:': [byte(240),159,136,178]
	':u7a7a:': [byte(240),159,136,179]
	':uganda:': [byte(240),159,135,186,240,159,135,172]
	':uk:': [byte(240),159,135,172,240,159,135,167]
	':ukraine:': [byte(240),159,135,186,240,159,135,166]
	':umbrella:': [byte(226),152,148]
	':unamused:': [byte(240),159,152,146]
	':underage:': [byte(240),159,148,158]
	':unicorn:': [byte(240),159,166,132]
	':united_arab_emirates:': [byte(240),159,135,166,240,159,135,170]
	':united_nations:': [byte(240),159,135,186,240,159,135,179]
	':unlock:': [byte(240),159,148,147]
	':up:': [byte(240),159,134,153]
	':upside_down_face:': [byte(240),159,153,131]
	':uruguay:': [byte(240),159,135,186,240,159,135,190]
	':us:': [byte(240),159,135,186,240,159,135,184]
	':us_outlying_islands:': [byte(240),159,135,186,240,159,135,178]
	':us_virgin_islands:': [byte(240),159,135,187,240,159,135,174]
	':uzbekistan:': [byte(240),159,135,186,240,159,135,191]
	':v:': [byte(226),156,140]
	':vampire:': [byte(240),159,167,155]
	':vampire_man:': [byte(240),159,167,155,226,153,130]
	':vampire_woman:': [byte(240),159,167,155,226,153,128]
	':vanuatu:': [byte(240),159,135,187,240,159,135,186]
	':vatican_city:': [byte(240),159,135,187,240,159,135,166]
	':venezuela:': [byte(240),159,135,187,240,159,135,170]
	':vertical_traffic_light:': [byte(240),159,154,166]
	':vhs:': [byte(240),159,147,188]
	':vibration_mode:': [byte(240),159,147,179]
	':video_camera:': [byte(240),159,147,185]
	':video_game:': [byte(240),159,142,174]
	':vietnam:': [byte(240),159,135,187,240,159,135,179]
	':violin:': [byte(240),159,142,187]
	':virgo:': [byte(226),153,141]
	':volcano:': [byte(240),159,140,139]
	':volleyball:': [byte(240),159,143,144]
	':vomiting_face:': [byte(240),159,164,174]
	':vs:': [byte(240),159,134,154]
	':vulcan_salute:': [byte(240),159,150,150]
	':waffle:': [byte(240),159,167,135]
	':wales:': [byte(240),159,143,180,243,160,129,167,243,160,129,162,243,160,129,183,243,160,129,172,243,160,129,179,243,160,129,191]
	':walking:': [byte(240),159,154,182]
	':walking_man:': [byte(240),159,154,182,226,153,130]
	':walking_woman:': [byte(240),159,154,182,226,153,128]
	':wallis_futuna:': [byte(240),159,135,188,240,159,135,171]
	':waning_crescent_moon:': [byte(240),159,140,152]
	':waning_gibbous_moon:': [byte(240),159,140,150]
	':warning:': [byte(226),154,160]
	':wastebasket:': [byte(240),159,151,145]
	':watch:': [byte(226),140,154]
	':water_buffalo:': [byte(240),159,144,131]
	':water_polo:': [byte(240),159,164,189]
	':watermelon:': [byte(240),159,141,137]
	':wave:': [byte(240),159,145,139]
	':wavy_dash:': [byte(227),128,176]
	':waxing_crescent_moon:': [byte(240),159,140,146]
	':waxing_gibbous_moon:': [byte(240),159,140,148]
	':wc:': [byte(240),159,154,190]
	':weary:': [byte(240),159,152,169]
	':wedding:': [byte(240),159,146,146]
	':weight_lifting:': [byte(240),159,143,139]
	':weight_lifting_man:': [byte(240),159,143,139,226,153,130]
	':weight_lifting_woman:': [byte(240),159,143,139,226,153,128]
	':western_sahara:': [byte(240),159,135,170,240,159,135,173]
	':whale:': [byte(240),159,144,179]
	':whale2:': [byte(240),159,144,139]
	':wheel_of_dharma:': [byte(226),152,184]
	':wheelchair:': [byte(226),153,191]
	':white_check_mark:': [byte(226),156,133]
	':white_circle:': [byte(226),154,170]
	':white_flag:': [byte(240),159,143,179]
	':white_flower:': [byte(240),159,146,174]
	':white_haired_man:': [byte(240),159,145,168,240,159,166,179]
	':white_haired_woman:': [byte(240),159,145,169,240,159,166,179]
	':white_heart:': [byte(240),159,164,141]
	':white_large_square:': [byte(226),172,156]
	':white_medium_small_square:': [byte(226),151,189]
	':white_medium_square:': [byte(226),151,187]
	':white_small_square:': [byte(226),150,171]
	':white_square_button:': [byte(240),159,148,179]
	':wilted_flower:': [byte(240),159,165,128]
	':wind_chime:': [byte(240),159,142,144]
	':wind_face:': [byte(240),159,140,172]
	':wine_glass:': [byte(240),159,141,183]
	':wink:': [byte(240),159,152,137]
	':wolf:': [byte(240),159,144,186]
	':woman:': [byte(240),159,145,169]
	':woman_artist:': [byte(240),159,145,169,240,159,142,168]
	':woman_astronaut:': [byte(240),159,145,169,240,159,154,128]
	':woman_cartwheeling:': [byte(240),159,164,184,226,153,128]
	':woman_cook:': [byte(240),159,145,169,240,159,141,179]
	':woman_dancing:': [byte(240),159,146,131]
	':woman_facepalming:': [byte(240),159,164,166,226,153,128]
	':woman_factory_worker:': [byte(240),159,145,169,240,159,143,173]
	':woman_farmer:': [byte(240),159,145,169,240,159,140,190]
	':woman_firefighter:': [byte(240),159,145,169,240,159,154,146]
	':woman_health_worker:': [byte(240),159,145,169,226,154,149]
	':woman_in_manual_wheelchair:': [byte(240),159,145,169,240,159,166,189]
	':woman_in_motorized_wheelchair:': [byte(240),159,145,169,240,159,166,188]
	':woman_judge:': [byte(240),159,145,169,226,154,150]
	':woman_juggling:': [byte(240),159,164,185,226,153,128]
	':woman_mechanic:': [byte(240),159,145,169,240,159,148,167]
	':woman_office_worker:': [byte(240),159,145,169,240,159,146,188]
	':woman_pilot:': [byte(240),159,145,169,226,156,136]
	':woman_playing_handball:': [byte(240),159,164,190,226,153,128]
	':woman_playing_water_polo:': [byte(240),159,164,189,226,153,128]
	':woman_scientist:': [byte(240),159,145,169,240,159,148,172]
	':woman_shrugging:': [byte(240),159,164,183,226,153,128]
	':woman_singer:': [byte(240),159,145,169,240,159,142,164]
	':woman_student:': [byte(240),159,145,169,240,159,142,147]
	':woman_teacher:': [byte(240),159,145,169,240,159,143,171]
	':woman_technologist:': [byte(240),159,145,169,240,159,146,187]
	':woman_with_headscarf:': [byte(240),159,167,149]
	':woman_with_probing_cane:': [byte(240),159,145,169,240,159,166,175]
	':woman_with_turban:': [byte(240),159,145,179,226,153,128]
	':womans_clothes:': [byte(240),159,145,154]
	':womans_hat:': [byte(240),159,145,146]
	':women_wrestling:': [byte(240),159,164,188,226,153,128]
	':womens:': [byte(240),159,154,186]
	':woozy_face:': [byte(240),159,165,180]
	':world_map:': [byte(240),159,151,186]
	':worried:': [byte(240),159,152,159]
	':wrench:': [byte(240),159,148,167]
	':wrestling:': [byte(240),159,164,188]
	':writing_hand:': [byte(226),156,141]
	':x:': [byte(226),157,140]
	':yarn:': [byte(240),159,167,182]
	':yawning_face:': [byte(240),159,165,177]
	':yellow_circle:': [byte(240),159,159,161]
	':yellow_heart:': [byte(240),159,146,155]
	':yellow_square:': [byte(240),159,159,168]
	':yemen:': [byte(240),159,135,190,240,159,135,170]
	':yen:': [byte(240),159,146,180]
	':yin_yang:': [byte(226),152,175]
	':yo_yo:': [byte(240),159,170,128]
	':yum:': [byte(240),159,152,139]
	':zambia:': [byte(240),159,135,191,240,159,135,178]
	':zany_face:': [byte(240),159,164,170]
	':zap:': [byte(226),154,161]
	':zebra:': [byte(240),159,166,147]
	':zero:': [byte(48),226,131,163]
	':zimbabwe:': [byte(240),159,135,191,240,159,135,188]
	':zipper_mouth_face:': [byte(240),159,164,144]
	':zombie:': [byte(240),159,167,159]
	':zombie_man:': [byte(240),159,167,159,226,153,130]
	':zombie_woman:': [byte(240),159,167,159,226,153,128]
	':zzz:': [byte(240),159,146,164]
}
