module moji

// https://api.github.com/emojis

pub const db = {
	'+1': '\xf0\x9f\x91\x8d',
	'-1': '\xf0\x9f\x91\x8e',
	'100': '\xf0\x9f\x92\xaf',
	'1234': '\xf0\x9f\x94\xa2',
	'1st_place_medal': '\xf0\x9f\xa5\x87',
	'2nd_place_medal': '\xf0\x9f\xa5\x88',
	'3rd_place_medal': '\xf0\x9f\xa5\x89',
	'8ball': '\xf0\x9f\x8e\xb1',
	'a': '\xf0\x9f\x85\xb0',
	'ab': '\xf0\x9f\x86\x8e',
	'abacus': '\xf0\x9f\xa7\xae',
	'abc': '\xf0\x9f\x94\xa4',
	'abcd': '\xf0\x9f\x94\xa1',
	'accept': '\xf0\x9f\x89\x91',
	'accordion': '\xf0\x9f\xaa\x97',
	'adhesive_bandage': '\xf0\x9f\xa9\xb9',
	'adult': '\xf0\x9f\xa7\x91',
	'aerial_tramway': '\xf0\x9f\x9a\xa1',
	'afghanistan': '\xf0\x9f\x87\xa6\xf0\x9f\x87\xab',
	'airplane': '\xe2\x9c\x88',
	'aland_islands': '\xf0\x9f\x87\xa6\xf0\x9f\x87\xbd',
	'alarm_clock': '\xe2\x8f\xb0',
	'albania': '\xf0\x9f\x87\xa6\xf0\x9f\x87\xb1',
	'alembic': '\xe2\x9a\x97',
	'algeria': '\xf0\x9f\x87\xa9\xf0\x9f\x87\xbf',
	'alien': '\xf0\x9f\x91\xbd',
	'ambulance': '\xf0\x9f\x9a\x91',
	'american_samoa': '\xf0\x9f\x87\xa6\xf0\x9f\x87\xb8',
	'amphora': '\xf0\x9f\x8f\xba',
	'anatomical_heart': '\xf0\x9f\xab\x80',
	'anchor': '\xe2\x9a\x93',
	'andorra': '\xf0\x9f\x87\xa6\xf0\x9f\x87\xa9',
	'angel': '\xf0\x9f\x91\xbc',
	'anger': '\xf0\x9f\x92\xa2',
	'angola': '\xf0\x9f\x87\xa6\xf0\x9f\x87\xb4',
	'angry': '\xf0\x9f\x98\xa0',
	'anguilla': '\xf0\x9f\x87\xa6\xf0\x9f\x87\xae',
	'anguished': '\xf0\x9f\x98\xa7',
	'ant': '\xf0\x9f\x90\x9c',
	'antarctica': '\xf0\x9f\x87\xa6\xf0\x9f\x87\xb6',
	'antigua_barbuda': '\xf0\x9f\x87\xa6\xf0\x9f\x87\xac',
	'apple': '\xf0\x9f\x8d\x8e',
	'aquarius': '\xe2\x99\x92',
	'argentina': '\xf0\x9f\x87\xa6\xf0\x9f\x87\xb7',
	'aries': '\xe2\x99\x88',
	'armenia': '\xf0\x9f\x87\xa6\xf0\x9f\x87\xb2',
	'arrow_backward': '\xe2\x97\x80',
	'arrow_double_down': '\xe2\x8f\xac',
	'arrow_double_up': '\xe2\x8f\xab',
	'arrow_down': '\xe2\xac\x87',
	'arrow_down_small': '\xf0\x9f\x94\xbd',
	'arrow_forward': '\xe2\x96\xb6',
	'arrow_heading_down': '\xe2\xa4\xb5',
	'arrow_heading_up': '\xe2\xa4\xb4',
	'arrow_left': '\xe2\xac\x85',
	'arrow_lower_left': '\xe2\x86\x99',
	'arrow_lower_right': '\xe2\x86\x98',
	'arrow_right': '\xe2\x9e\xa1',
	'arrow_right_hook': '\xe2\x86\xaa',
	'arrow_up': '\xe2\xac\x86',
	'arrow_up_down': '\xe2\x86\x95',
	'arrow_up_small': '\xf0\x9f\x94\xbc',
	'arrow_upper_left': '\xe2\x86\x96',
	'arrow_upper_right': '\xe2\x86\x97',
	'arrows_clockwise': '\xf0\x9f\x94\x83',
	'arrows_counterclockwise': '\xf0\x9f\x94\x84',
	'art': '\xf0\x9f\x8e\xa8',
	'articulated_lorry': '\xf0\x9f\x9a\x9b',
	'artificial_satellite': '\xf0\x9f\x9b\xb0',
	'artist': '\xf0\x9f\xa7\x91\xf0\x9f\x8e\xa8',
	'aruba': '\xf0\x9f\x87\xa6\xf0\x9f\x87\xbc',
	'ascension_island': '\xf0\x9f\x87\xa6\xf0\x9f\x87\xa8',
	'asterisk': '\x2a\xe2\x83\xa3',
	'astonished': '\xf0\x9f\x98\xb2',
	'astronaut': '\xf0\x9f\xa7\x91\xf0\x9f\x9a\x80',
	'athletic_shoe': '\xf0\x9f\x91\x9f',
	'atm': '\xf0\x9f\x8f\xa7',
	'atom_symbol': '\xe2\x9a\x9b',
	'australia': '\xf0\x9f\x87\xa6\xf0\x9f\x87\xba',
	'austria': '\xf0\x9f\x87\xa6\xf0\x9f\x87\xb9',
	'auto_rickshaw': '\xf0\x9f\x9b\xba',
	'avocado': '\xf0\x9f\xa5\x91',
	'axe': '\xf0\x9f\xaa\x93',
	'azerbaijan': '\xf0\x9f\x87\xa6\xf0\x9f\x87\xbf',
	'b': '\xf0\x9f\x85\xb1',
	'baby': '\xf0\x9f\x91\xb6',
	'baby_bottle': '\xf0\x9f\x8d\xbc',
	'baby_chick': '\xf0\x9f\x90\xa4',
	'baby_symbol': '\xf0\x9f\x9a\xbc',
	'back': '\xf0\x9f\x94\x99',
	'bacon': '\xf0\x9f\xa5\x93',
	'badger': '\xf0\x9f\xa6\xa1',
	'badminton': '\xf0\x9f\x8f\xb8',
	'bagel': '\xf0\x9f\xa5\xaf',
	'baggage_claim': '\xf0\x9f\x9b\x84',
	'baguette_bread': '\xf0\x9f\xa5\x96',
	'bahamas': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xb8',
	'bahrain': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xad',
	'balance_scale': '\xe2\x9a\x96',
	'bald_man': '\xf0\x9f\x91\xa8\xf0\x9f\xa6\xb2',
	'bald_woman': '\xf0\x9f\x91\xa9\xf0\x9f\xa6\xb2',
	'ballet_shoes': '\xf0\x9f\xa9\xb0',
	'balloon': '\xf0\x9f\x8e\x88',
	'ballot_box': '\xf0\x9f\x97\xb3',
	'ballot_box_with_check': '\xe2\x98\x91',
	'bamboo': '\xf0\x9f\x8e\x8d',
	'banana': '\xf0\x9f\x8d\x8c',
	'bangbang': '\xe2\x80\xbc',
	'bangladesh': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xa9',
	'banjo': '\xf0\x9f\xaa\x95',
	'bank': '\xf0\x9f\x8f\xa6',
	'bar_chart': '\xf0\x9f\x93\x8a',
	'barbados': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xa7',
	'barber': '\xf0\x9f\x92\x88',
	'baseball': '\xe2\x9a\xbe',
	'basket': '\xf0\x9f\xa7\xba',
	'basketball': '\xf0\x9f\x8f\x80',
	'basketball_man': '\xe2\x9b\xb9\xe2\x99\x82',
	'basketball_woman': '\xe2\x9b\xb9\xe2\x99\x80',
	'bat': '\xf0\x9f\xa6\x87',
	'bath': '\xf0\x9f\x9b\x80',
	'bathtub': '\xf0\x9f\x9b\x81',
	'battery': '\xf0\x9f\x94\x8b',
	'beach_umbrella': '\xf0\x9f\x8f\x96',
	'bear': '\xf0\x9f\x90\xbb',
	'bearded_person': '\xf0\x9f\xa7\x94',
	'beaver': '\xf0\x9f\xa6\xab',
	'bed': '\xf0\x9f\x9b\x8f',
	'bee': '\xf0\x9f\x90\x9d',
	'beer': '\xf0\x9f\x8d\xba',
	'beers': '\xf0\x9f\x8d\xbb',
	'beetle': '\xf0\x9f\xaa\xb2',
	'beginner': '\xf0\x9f\x94\xb0',
	'belarus': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xbe',
	'belgium': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xaa',
	'belize': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xbf',
	'bell': '\xf0\x9f\x94\x94',
	'bell_pepper': '\xf0\x9f\xab\x91',
	'bellhop_bell': '\xf0\x9f\x9b\x8e',
	'benin': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xaf',
	'bento': '\xf0\x9f\x8d\xb1',
	'bermuda': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xb2',
	'beverage_box': '\xf0\x9f\xa7\x83',
	'bhutan': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xb9',
	'bicyclist': '\xf0\x9f\x9a\xb4',
	'bike': '\xf0\x9f\x9a\xb2',
	'biking_man': '\xf0\x9f\x9a\xb4\xe2\x99\x82',
	'biking_woman': '\xf0\x9f\x9a\xb4\xe2\x99\x80',
	'bikini': '\xf0\x9f\x91\x99',
	'billed_cap': '\xf0\x9f\xa7\xa2',
	'biohazard': '\xe2\x98\xa3',
	'bird': '\xf0\x9f\x90\xa6',
	'birthday': '\xf0\x9f\x8e\x82',
	'bison': '\xf0\x9f\xa6\xac',
	'black_cat': '\xf0\x9f\x90\x88\xe2\xac\x9b',
	'black_circle': '\xe2\x9a\xab',
	'black_flag': '\xf0\x9f\x8f\xb4',
	'black_heart': '\xf0\x9f\x96\xa4',
	'black_joker': '\xf0\x9f\x83\x8f',
	'black_large_square': '\xe2\xac\x9b',
	'black_medium_small_square': '\xe2\x97\xbe',
	'black_medium_square': '\xe2\x97\xbc',
	'black_nib': '\xe2\x9c\x92',
	'black_small_square': '\xe2\x96\xaa',
	'black_square_button': '\xf0\x9f\x94\xb2',
	'blond_haired_man': '\xf0\x9f\x91\xb1\xe2\x99\x82',
	'blond_haired_person': '\xf0\x9f\x91\xb1',
	'blond_haired_woman': '\xf0\x9f\x91\xb1\xe2\x99\x80',
	'blonde_woman': '\xf0\x9f\x91\xb1\xe2\x99\x80',
	'blossom': '\xf0\x9f\x8c\xbc',
	'blowfish': '\xf0\x9f\x90\xa1',
	'blue_book': '\xf0\x9f\x93\x98',
	'blue_car': '\xf0\x9f\x9a\x99',
	'blue_heart': '\xf0\x9f\x92\x99',
	'blue_square': '\xf0\x9f\x9f\xa6',
	'blueberries': '\xf0\x9f\xab\x90',
	'blush': '\xf0\x9f\x98\x8a',
	'boar': '\xf0\x9f\x90\x97',
	'boat': '\xe2\x9b\xb5',
	'bolivia': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xb4',
	'bomb': '\xf0\x9f\x92\xa3',
	'bone': '\xf0\x9f\xa6\xb4',
	'book': '\xf0\x9f\x93\x96',
	'bookmark': '\xf0\x9f\x94\x96',
	'bookmark_tabs': '\xf0\x9f\x93\x91',
	'books': '\xf0\x9f\x93\x9a',
	'boom': '\xf0\x9f\x92\xa5',
	'boomerang': '\xf0\x9f\xaa\x83',
	'boot': '\xf0\x9f\x91\xa2',
	'bosnia_herzegovina': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xa6',
	'botswana': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xbc',
	'bouncing_ball_man': '\xe2\x9b\xb9\xe2\x99\x82',
	'bouncing_ball_person': '\xe2\x9b\xb9',
	'bouncing_ball_woman': '\xe2\x9b\xb9\xe2\x99\x80',
	'bouquet': '\xf0\x9f\x92\x90',
	'bouvet_island': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xbb',
	'bow': '\xf0\x9f\x99\x87',
	'bow_and_arrow': '\xf0\x9f\x8f\xb9',
	'bowing_man': '\xf0\x9f\x99\x87\xe2\x99\x82',
	'bowing_woman': '\xf0\x9f\x99\x87\xe2\x99\x80',
	'bowl_with_spoon': '\xf0\x9f\xa5\xa3',
	'bowling': '\xf0\x9f\x8e\xb3',
	'boxing_glove': '\xf0\x9f\xa5\x8a',
	'boy': '\xf0\x9f\x91\xa6',
	'brain': '\xf0\x9f\xa7\xa0',
	'brazil': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xb7',
	'bread': '\xf0\x9f\x8d\x9e',
	'breast_feeding': '\xf0\x9f\xa4\xb1',
	'bricks': '\xf0\x9f\xa7\xb1',
	'bride_with_veil': '\xf0\x9f\x91\xb0\xe2\x99\x80',
	'bridge_at_night': '\xf0\x9f\x8c\x89',
	'briefcase': '\xf0\x9f\x92\xbc',
	'british_indian_ocean_territory': '\xf0\x9f\x87\xae\xf0\x9f\x87\xb4',
	'british_virgin_islands': '\xf0\x9f\x87\xbb\xf0\x9f\x87\xac',
	'broccoli': '\xf0\x9f\xa5\xa6',
	'broken_heart': '\xf0\x9f\x92\x94',
	'broom': '\xf0\x9f\xa7\xb9',
	'brown_circle': '\xf0\x9f\x9f\xa4',
	'brown_heart': '\xf0\x9f\xa4\x8e',
	'brown_square': '\xf0\x9f\x9f\xab',
	'brunei': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xb3',
	'bubble_tea': '\xf0\x9f\xa7\x8b',
	'bucket': '\xf0\x9f\xaa\xa3',
	'bug': '\xf0\x9f\x90\x9b',
	'building_construction': '\xf0\x9f\x8f\x97',
	'bulb': '\xf0\x9f\x92\xa1',
	'bulgaria': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xac',
	'bullettrain_front': '\xf0\x9f\x9a\x85',
	'bullettrain_side': '\xf0\x9f\x9a\x84',
	'burkina_faso': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xab',
	'burrito': '\xf0\x9f\x8c\xaf',
	'burundi': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xae',
	'bus': '\xf0\x9f\x9a\x8c',
	'business_suit_levitating': '\xf0\x9f\x95\xb4',
	'busstop': '\xf0\x9f\x9a\x8f',
	'bust_in_silhouette': '\xf0\x9f\x91\xa4',
	'busts_in_silhouette': '\xf0\x9f\x91\xa5',
	'butter': '\xf0\x9f\xa7\x88',
	'butterfly': '\xf0\x9f\xa6\x8b',
	'cactus': '\xf0\x9f\x8c\xb5',
	'cake': '\xf0\x9f\x8d\xb0',
	'calendar': '\xf0\x9f\x93\x86',
	'call_me_hand': '\xf0\x9f\xa4\x99',
	'calling': '\xf0\x9f\x93\xb2',
	'cambodia': '\xf0\x9f\x87\xb0\xf0\x9f\x87\xad',
	'camel': '\xf0\x9f\x90\xab',
	'camera': '\xf0\x9f\x93\xb7',
	'camera_flash': '\xf0\x9f\x93\xb8',
	'cameroon': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xb2',
	'camping': '\xf0\x9f\x8f\x95',
	'canada': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xa6',
	'canary_islands': '\xf0\x9f\x87\xae\xf0\x9f\x87\xa8',
	'cancer': '\xe2\x99\x8b',
	'candle': '\xf0\x9f\x95\xaf',
	'candy': '\xf0\x9f\x8d\xac',
	'canned_food': '\xf0\x9f\xa5\xab',
	'canoe': '\xf0\x9f\x9b\xb6',
	'cape_verde': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xbb',
	'capital_abcd': '\xf0\x9f\x94\xa0',
	'capricorn': '\xe2\x99\x91',
	'car': '\xf0\x9f\x9a\x97',
	'card_file_box': '\xf0\x9f\x97\x83',
	'card_index': '\xf0\x9f\x93\x87',
	'card_index_dividers': '\xf0\x9f\x97\x82',
	'caribbean_netherlands': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xb6',
	'carousel_horse': '\xf0\x9f\x8e\xa0',
	'carpentry_saw': '\xf0\x9f\xaa\x9a',
	'carrot': '\xf0\x9f\xa5\x95',
	'cartwheeling': '\xf0\x9f\xa4\xb8',
	'cat': '\xf0\x9f\x90\xb1',
	'cat2': '\xf0\x9f\x90\x88',
	'cayman_islands': '\xf0\x9f\x87\xb0\xf0\x9f\x87\xbe',
	'cd': '\xf0\x9f\x92\xbf',
	'central_african_republic': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xab',
	'ceuta_melilla': '\xf0\x9f\x87\xaa\xf0\x9f\x87\xa6',
	'chad': '\xf0\x9f\x87\xb9\xf0\x9f\x87\xa9',
	'chains': '\xe2\x9b\x93',
	'chair': '\xf0\x9f\xaa\x91',
	'champagne': '\xf0\x9f\x8d\xbe',
	'chart': '\xf0\x9f\x92\xb9',
	'chart_with_downwards_trend': '\xf0\x9f\x93\x89',
	'chart_with_upwards_trend': '\xf0\x9f\x93\x88',
	'checkered_flag': '\xf0\x9f\x8f\x81',
	'cheese': '\xf0\x9f\xa7\x80',
	'cherries': '\xf0\x9f\x8d\x92',
	'cherry_blossom': '\xf0\x9f\x8c\xb8',
	'chess_pawn': '\xe2\x99\x9f',
	'chestnut': '\xf0\x9f\x8c\xb0',
	'chicken': '\xf0\x9f\x90\x94',
	'child': '\xf0\x9f\xa7\x92',
	'children_crossing': '\xf0\x9f\x9a\xb8',
	'chile': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xb1',
	'chipmunk': '\xf0\x9f\x90\xbf',
	'chocolate_bar': '\xf0\x9f\x8d\xab',
	'chopsticks': '\xf0\x9f\xa5\xa2',
	'christmas_island': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xbd',
	'christmas_tree': '\xf0\x9f\x8e\x84',
	'church': '\xe2\x9b\xaa',
	'cinema': '\xf0\x9f\x8e\xa6',
	'circus_tent': '\xf0\x9f\x8e\xaa',
	'city_sunrise': '\xf0\x9f\x8c\x87',
	'city_sunset': '\xf0\x9f\x8c\x86',
	'cityscape': '\xf0\x9f\x8f\x99',
	'cl': '\xf0\x9f\x86\x91',
	'clamp': '\xf0\x9f\x97\x9c',
	'clap': '\xf0\x9f\x91\x8f',
	'clapper': '\xf0\x9f\x8e\xac',
	'classical_building': '\xf0\x9f\x8f\x9b',
	'climbing': '\xf0\x9f\xa7\x97',
	'climbing_man': '\xf0\x9f\xa7\x97\xe2\x99\x82',
	'climbing_woman': '\xf0\x9f\xa7\x97\xe2\x99\x80',
	'clinking_glasses': '\xf0\x9f\xa5\x82',
	'clipboard': '\xf0\x9f\x93\x8b',
	'clipperton_island': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xb5',
	'clock1': '\xf0\x9f\x95\x90',
	'clock10': '\xf0\x9f\x95\x99',
	'clock1030': '\xf0\x9f\x95\xa5',
	'clock11': '\xf0\x9f\x95\x9a',
	'clock1130': '\xf0\x9f\x95\xa6',
	'clock12': '\xf0\x9f\x95\x9b',
	'clock1230': '\xf0\x9f\x95\xa7',
	'clock130': '\xf0\x9f\x95\x9c',
	'clock2': '\xf0\x9f\x95\x91',
	'clock230': '\xf0\x9f\x95\x9d',
	'clock3': '\xf0\x9f\x95\x92',
	'clock330': '\xf0\x9f\x95\x9e',
	'clock4': '\xf0\x9f\x95\x93',
	'clock430': '\xf0\x9f\x95\x9f',
	'clock5': '\xf0\x9f\x95\x94',
	'clock530': '\xf0\x9f\x95\xa0',
	'clock6': '\xf0\x9f\x95\x95',
	'clock630': '\xf0\x9f\x95\xa1',
	'clock7': '\xf0\x9f\x95\x96',
	'clock730': '\xf0\x9f\x95\xa2',
	'clock8': '\xf0\x9f\x95\x97',
	'clock830': '\xf0\x9f\x95\xa3',
	'clock9': '\xf0\x9f\x95\x98',
	'clock930': '\xf0\x9f\x95\xa4',
	'closed_book': '\xf0\x9f\x93\x95',
	'closed_lock_with_key': '\xf0\x9f\x94\x90',
	'closed_umbrella': '\xf0\x9f\x8c\x82',
	'cloud': '\xe2\x98\x81',
	'cloud_with_lightning': '\xf0\x9f\x8c\xa9',
	'cloud_with_lightning_and_rain': '\xe2\x9b\x88',
	'cloud_with_rain': '\xf0\x9f\x8c\xa7',
	'cloud_with_snow': '\xf0\x9f\x8c\xa8',
	'clown_face': '\xf0\x9f\xa4\xa1',
	'clubs': '\xe2\x99\xa3',
	'cn': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xb3',
	'coat': '\xf0\x9f\xa7\xa5',
	'cockroach': '\xf0\x9f\xaa\xb3',
	'cocktail': '\xf0\x9f\x8d\xb8',
	'coconut': '\xf0\x9f\xa5\xa5',
	'cocos_islands': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xa8',
	'coffee': '\xe2\x98\x95',
	'coffin': '\xe2\x9a\xb0',
	'coin': '\xf0\x9f\xaa\x99',
	'cold_face': '\xf0\x9f\xa5\xb6',
	'cold_sweat': '\xf0\x9f\x98\xb0',
	'collision': '\xf0\x9f\x92\xa5',
	'colombia': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xb4',
	'comet': '\xe2\x98\x84',
	'comoros': '\xf0\x9f\x87\xb0\xf0\x9f\x87\xb2',
	'compass': '\xf0\x9f\xa7\xad',
	'computer': '\xf0\x9f\x92\xbb',
	'computer_mouse': '\xf0\x9f\x96\xb1',
	'confetti_ball': '\xf0\x9f\x8e\x8a',
	'confounded': '\xf0\x9f\x98\x96',
	'confused': '\xf0\x9f\x98\x95',
	'congo_brazzaville': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xac',
	'congo_kinshasa': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xa9',
	'congratulations': '\xe3\x8a\x97',
	'construction': '\xf0\x9f\x9a\xa7',
	'construction_worker': '\xf0\x9f\x91\xb7',
	'construction_worker_man': '\xf0\x9f\x91\xb7\xe2\x99\x82',
	'construction_worker_woman': '\xf0\x9f\x91\xb7\xe2\x99\x80',
	'control_knobs': '\xf0\x9f\x8e\x9b',
	'convenience_store': '\xf0\x9f\x8f\xaa',
	'cook': '\xf0\x9f\xa7\x91\xf0\x9f\x8d\xb3',
	'cook_islands': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xb0',
	'cookie': '\xf0\x9f\x8d\xaa',
	'cool': '\xf0\x9f\x86\x92',
	'cop': '\xf0\x9f\x91\xae',
	'copyright': '\xc2\xa9',
	'corn': '\xf0\x9f\x8c\xbd',
	'costa_rica': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xb7',
	'cote_divoire': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xae',
	'couch_and_lamp': '\xf0\x9f\x9b\x8b',
	'couple': '\xf0\x9f\x91\xab',
	'couple_with_heart': '\xf0\x9f\x92\x91',
	'couple_with_heart_man_man': '\xf0\x9f\x91\xa8\xe2\x9d\xa4\xf0\x9f\x91\xa8',
	'couple_with_heart_woman_man': '\xf0\x9f\x91\xa9\xe2\x9d\xa4\xf0\x9f\x91\xa8',
	'couple_with_heart_woman_woman': '\xf0\x9f\x91\xa9\xe2\x9d\xa4\xf0\x9f\x91\xa9',
	'couplekiss': '\xf0\x9f\x92\x8f',
	'couplekiss_man_man': '\xf0\x9f\x91\xa8\xe2\x9d\xa4\xf0\x9f\x92\x8b\xf0\x9f\x91\xa8',
	'couplekiss_man_woman': '\xf0\x9f\x91\xa9\xe2\x9d\xa4\xf0\x9f\x92\x8b\xf0\x9f\x91\xa8',
	'couplekiss_woman_woman': '\xf0\x9f\x91\xa9\xe2\x9d\xa4\xf0\x9f\x92\x8b\xf0\x9f\x91\xa9',
	'cow': '\xf0\x9f\x90\xae',
	'cow2': '\xf0\x9f\x90\x84',
	'cowboy_hat_face': '\xf0\x9f\xa4\xa0',
	'crab': '\xf0\x9f\xa6\x80',
	'crayon': '\xf0\x9f\x96\x8d',
	'credit_card': '\xf0\x9f\x92\xb3',
	'crescent_moon': '\xf0\x9f\x8c\x99',
	'cricket': '\xf0\x9f\xa6\x97',
	'cricket_game': '\xf0\x9f\x8f\x8f',
	'croatia': '\xf0\x9f\x87\xad\xf0\x9f\x87\xb7',
	'crocodile': '\xf0\x9f\x90\x8a',
	'croissant': '\xf0\x9f\xa5\x90',
	'crossed_fingers': '\xf0\x9f\xa4\x9e',
	'crossed_flags': '\xf0\x9f\x8e\x8c',
	'crossed_swords': '\xe2\x9a\x94',
	'crown': '\xf0\x9f\x91\x91',
	'cry': '\xf0\x9f\x98\xa2',
	'crying_cat_face': '\xf0\x9f\x98\xbf',
	'crystal_ball': '\xf0\x9f\x94\xae',
	'cuba': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xba',
	'cucumber': '\xf0\x9f\xa5\x92',
	'cup_with_straw': '\xf0\x9f\xa5\xa4',
	'cupcake': '\xf0\x9f\xa7\x81',
	'cupid': '\xf0\x9f\x92\x98',
	'curacao': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xbc',
	'curling_stone': '\xf0\x9f\xa5\x8c',
	'curly_haired_man': '\xf0\x9f\x91\xa8\xf0\x9f\xa6\xb1',
	'curly_haired_woman': '\xf0\x9f\x91\xa9\xf0\x9f\xa6\xb1',
	'curly_loop': '\xe2\x9e\xb0',
	'currency_exchange': '\xf0\x9f\x92\xb1',
	'curry': '\xf0\x9f\x8d\x9b',
	'cursing_face': '\xf0\x9f\xa4\xac',
	'custard': '\xf0\x9f\x8d\xae',
	'customs': '\xf0\x9f\x9b\x83',
	'cut_of_meat': '\xf0\x9f\xa5\xa9',
	'cyclone': '\xf0\x9f\x8c\x80',
	'cyprus': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xbe',
	'czech_republic': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xbf',
	'dagger': '\xf0\x9f\x97\xa1',
	'dancer': '\xf0\x9f\x92\x83',
	'dancers': '\xf0\x9f\x91\xaf',
	'dancing_men': '\xf0\x9f\x91\xaf\xe2\x99\x82',
	'dancing_women': '\xf0\x9f\x91\xaf\xe2\x99\x80',
	'dango': '\xf0\x9f\x8d\xa1',
	'dark_sunglasses': '\xf0\x9f\x95\xb6',
	'dart': '\xf0\x9f\x8e\xaf',
	'dash': '\xf0\x9f\x92\xa8',
	'date': '\xf0\x9f\x93\x85',
	'de': '\xf0\x9f\x87\xa9\xf0\x9f\x87\xaa',
	'deaf_man': '\xf0\x9f\xa7\x8f\xe2\x99\x82',
	'deaf_person': '\xf0\x9f\xa7\x8f',
	'deaf_woman': '\xf0\x9f\xa7\x8f\xe2\x99\x80',
	'deciduous_tree': '\xf0\x9f\x8c\xb3',
	'deer': '\xf0\x9f\xa6\x8c',
	'denmark': '\xf0\x9f\x87\xa9\xf0\x9f\x87\xb0',
	'department_store': '\xf0\x9f\x8f\xac',
	'derelict_house': '\xf0\x9f\x8f\x9a',
	'desert': '\xf0\x9f\x8f\x9c',
	'desert_island': '\xf0\x9f\x8f\x9d',
	'desktop_computer': '\xf0\x9f\x96\xa5',
	'detective': '\xf0\x9f\x95\xb5',
	'diamond_shape_with_a_dot_inside': '\xf0\x9f\x92\xa0',
	'diamonds': '\xe2\x99\xa6',
	'diego_garcia': '\xf0\x9f\x87\xa9\xf0\x9f\x87\xac',
	'disappointed': '\xf0\x9f\x98\x9e',
	'disappointed_relieved': '\xf0\x9f\x98\xa5',
	'disguised_face': '\xf0\x9f\xa5\xb8',
	'diving_mask': '\xf0\x9f\xa4\xbf',
	'diya_lamp': '\xf0\x9f\xaa\x94',
	'dizzy': '\xf0\x9f\x92\xab',
	'dizzy_face': '\xf0\x9f\x98\xb5',
	'djibouti': '\xf0\x9f\x87\xa9\xf0\x9f\x87\xaf',
	'dna': '\xf0\x9f\xa7\xac',
	'do_not_litter': '\xf0\x9f\x9a\xaf',
	'dodo': '\xf0\x9f\xa6\xa4',
	'dog': '\xf0\x9f\x90\xb6',
	'dog2': '\xf0\x9f\x90\x95',
	'dollar': '\xf0\x9f\x92\xb5',
	'dolls': '\xf0\x9f\x8e\x8e',
	'dolphin': '\xf0\x9f\x90\xac',
	'dominica': '\xf0\x9f\x87\xa9\xf0\x9f\x87\xb2',
	'dominican_republic': '\xf0\x9f\x87\xa9\xf0\x9f\x87\xb4',
	'door': '\xf0\x9f\x9a\xaa',
	'doughnut': '\xf0\x9f\x8d\xa9',
	'dove': '\xf0\x9f\x95\x8a',
	'dragon': '\xf0\x9f\x90\x89',
	'dragon_face': '\xf0\x9f\x90\xb2',
	'dress': '\xf0\x9f\x91\x97',
	'dromedary_camel': '\xf0\x9f\x90\xaa',
	'drooling_face': '\xf0\x9f\xa4\xa4',
	'drop_of_blood': '\xf0\x9f\xa9\xb8',
	'droplet': '\xf0\x9f\x92\xa7',
	'drum': '\xf0\x9f\xa5\x81',
	'duck': '\xf0\x9f\xa6\x86',
	'dumpling': '\xf0\x9f\xa5\x9f',
	'dvd': '\xf0\x9f\x93\x80',
	'e-mail': '\xf0\x9f\x93\xa7',
	'eagle': '\xf0\x9f\xa6\x85',
	'ear': '\xf0\x9f\x91\x82',
	'ear_of_rice': '\xf0\x9f\x8c\xbe',
	'ear_with_hearing_aid': '\xf0\x9f\xa6\xbb',
	'earth_africa': '\xf0\x9f\x8c\x8d',
	'earth_americas': '\xf0\x9f\x8c\x8e',
	'earth_asia': '\xf0\x9f\x8c\x8f',
	'ecuador': '\xf0\x9f\x87\xaa\xf0\x9f\x87\xa8',
	'egg': '\xf0\x9f\xa5\x9a',
	'eggplant': '\xf0\x9f\x8d\x86',
	'egypt': '\xf0\x9f\x87\xaa\xf0\x9f\x87\xac',
	'eight': '\x38\xe2\x83\xa3',
	'eight_pointed_black_star': '\xe2\x9c\xb4',
	'eight_spoked_asterisk': '\xe2\x9c\xb3',
	'eject_button': '\xe2\x8f\x8f',
	'el_salvador': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xbb',
	'electric_plug': '\xf0\x9f\x94\x8c',
	'elephant': '\xf0\x9f\x90\x98',
	'elevator': '\xf0\x9f\x9b\x97',
	'elf': '\xf0\x9f\xa7\x9d',
	'elf_man': '\xf0\x9f\xa7\x9d\xe2\x99\x82',
	'elf_woman': '\xf0\x9f\xa7\x9d\xe2\x99\x80',
	'email': '\xf0\x9f\x93\xa7',
	'end': '\xf0\x9f\x94\x9a',
	'england': '\xf0\x9f\x8f\xb4\xf3\xa0\x81\xa7\xf3\xa0\x81\xa2\xf3\xa0\x81\xa5\xf3\xa0\x81\xae\xf3\xa0\x81\xa7\xf3\xa0\x81\xbf',
	'envelope': '\xe2\x9c\x89',
	'envelope_with_arrow': '\xf0\x9f\x93\xa9',
	'equatorial_guinea': '\xf0\x9f\x87\xac\xf0\x9f\x87\xb6',
	'eritrea': '\xf0\x9f\x87\xaa\xf0\x9f\x87\xb7',
	'es': '\xf0\x9f\x87\xaa\xf0\x9f\x87\xb8',
	'estonia': '\xf0\x9f\x87\xaa\xf0\x9f\x87\xaa',
	'ethiopia': '\xf0\x9f\x87\xaa\xf0\x9f\x87\xb9',
	'eu': '\xf0\x9f\x87\xaa\xf0\x9f\x87\xba',
	'euro': '\xf0\x9f\x92\xb6',
	'european_castle': '\xf0\x9f\x8f\xb0',
	'european_post_office': '\xf0\x9f\x8f\xa4',
	'european_union': '\xf0\x9f\x87\xaa\xf0\x9f\x87\xba',
	'evergreen_tree': '\xf0\x9f\x8c\xb2',
	'exclamation': '\xe2\x9d\x97',
	'exploding_head': '\xf0\x9f\xa4\xaf',
	'expressionless': '\xf0\x9f\x98\x91',
	'eye': '\xf0\x9f\x91\x81',
	'eye_speech_bubble': '\xf0\x9f\x91\x81\xf0\x9f\x97\xa8',
	'eyeglasses': '\xf0\x9f\x91\x93',
	'eyes': '\xf0\x9f\x91\x80',
	'face_exhaling': '\xf0\x9f\x98\xae\xf0\x9f\x92\xa8',
	'face_in_clouds': '\xf0\x9f\x98\xb6\xf0\x9f\x8c\xab',
	'face_with_head_bandage': '\xf0\x9f\xa4\x95',
	'face_with_spiral_eyes': '\xf0\x9f\x98\xb5\xf0\x9f\x92\xab',
	'face_with_thermometer': '\xf0\x9f\xa4\x92',
	'facepalm': '\xf0\x9f\xa4\xa6',
	'facepunch': '\xf0\x9f\x91\x8a',
	'factory': '\xf0\x9f\x8f\xad',
	'factory_worker': '\xf0\x9f\xa7\x91\xf0\x9f\x8f\xad',
	'fairy': '\xf0\x9f\xa7\x9a',
	'fairy_man': '\xf0\x9f\xa7\x9a\xe2\x99\x82',
	'fairy_woman': '\xf0\x9f\xa7\x9a\xe2\x99\x80',
	'falafel': '\xf0\x9f\xa7\x86',
	'falkland_islands': '\xf0\x9f\x87\xab\xf0\x9f\x87\xb0',
	'fallen_leaf': '\xf0\x9f\x8d\x82',
	'family': '\xf0\x9f\x91\xaa',
	'family_man_boy': '\xf0\x9f\x91\xa8\xf0\x9f\x91\xa6',
	'family_man_boy_boy': '\xf0\x9f\x91\xa8\xf0\x9f\x91\xa6\xf0\x9f\x91\xa6',
	'family_man_girl': '\xf0\x9f\x91\xa8\xf0\x9f\x91\xa7',
	'family_man_girl_boy': '\xf0\x9f\x91\xa8\xf0\x9f\x91\xa7\xf0\x9f\x91\xa6',
	'family_man_girl_girl': '\xf0\x9f\x91\xa8\xf0\x9f\x91\xa7\xf0\x9f\x91\xa7',
	'family_man_man_boy': '\xf0\x9f\x91\xa8\xf0\x9f\x91\xa8\xf0\x9f\x91\xa6',
	'family_man_man_boy_boy': '\xf0\x9f\x91\xa8\xf0\x9f\x91\xa8\xf0\x9f\x91\xa6\xf0\x9f\x91\xa6',
	'family_man_man_girl': '\xf0\x9f\x91\xa8\xf0\x9f\x91\xa8\xf0\x9f\x91\xa7',
	'family_man_man_girl_boy': '\xf0\x9f\x91\xa8\xf0\x9f\x91\xa8\xf0\x9f\x91\xa7\xf0\x9f\x91\xa6',
	'family_man_man_girl_girl': '\xf0\x9f\x91\xa8\xf0\x9f\x91\xa8\xf0\x9f\x91\xa7\xf0\x9f\x91\xa7',
	'family_man_woman_boy': '\xf0\x9f\x91\xa8\xf0\x9f\x91\xa9\xf0\x9f\x91\xa6',
	'family_man_woman_boy_boy': '\xf0\x9f\x91\xa8\xf0\x9f\x91\xa9\xf0\x9f\x91\xa6\xf0\x9f\x91\xa6',
	'family_man_woman_girl': '\xf0\x9f\x91\xa8\xf0\x9f\x91\xa9\xf0\x9f\x91\xa7',
	'family_man_woman_girl_boy': '\xf0\x9f\x91\xa8\xf0\x9f\x91\xa9\xf0\x9f\x91\xa7\xf0\x9f\x91\xa6',
	'family_man_woman_girl_girl': '\xf0\x9f\x91\xa8\xf0\x9f\x91\xa9\xf0\x9f\x91\xa7\xf0\x9f\x91\xa7',
	'family_woman_boy': '\xf0\x9f\x91\xa9\xf0\x9f\x91\xa6',
	'family_woman_boy_boy': '\xf0\x9f\x91\xa9\xf0\x9f\x91\xa6\xf0\x9f\x91\xa6',
	'family_woman_girl': '\xf0\x9f\x91\xa9\xf0\x9f\x91\xa7',
	'family_woman_girl_boy': '\xf0\x9f\x91\xa9\xf0\x9f\x91\xa7\xf0\x9f\x91\xa6',
	'family_woman_girl_girl': '\xf0\x9f\x91\xa9\xf0\x9f\x91\xa7\xf0\x9f\x91\xa7',
	'family_woman_woman_boy': '\xf0\x9f\x91\xa9\xf0\x9f\x91\xa9\xf0\x9f\x91\xa6',
	'family_woman_woman_boy_boy': '\xf0\x9f\x91\xa9\xf0\x9f\x91\xa9\xf0\x9f\x91\xa6\xf0\x9f\x91\xa6',
	'family_woman_woman_girl': '\xf0\x9f\x91\xa9\xf0\x9f\x91\xa9\xf0\x9f\x91\xa7',
	'family_woman_woman_girl_boy': '\xf0\x9f\x91\xa9\xf0\x9f\x91\xa9\xf0\x9f\x91\xa7\xf0\x9f\x91\xa6',
	'family_woman_woman_girl_girl': '\xf0\x9f\x91\xa9\xf0\x9f\x91\xa9\xf0\x9f\x91\xa7\xf0\x9f\x91\xa7',
	'farmer': '\xf0\x9f\xa7\x91\xf0\x9f\x8c\xbe',
	'faroe_islands': '\xf0\x9f\x87\xab\xf0\x9f\x87\xb4',
	'fast_forward': '\xe2\x8f\xa9',
	'fax': '\xf0\x9f\x93\xa0',
	'fearful': '\xf0\x9f\x98\xa8',
	'feather': '\xf0\x9f\xaa\xb6',
	'feet': '\xf0\x9f\x90\xbe',
	'female_detective': '\xf0\x9f\x95\xb5\xe2\x99\x80',
	'female_sign': '\xe2\x99\x80',
	'ferris_wheel': '\xf0\x9f\x8e\xa1',
	'ferry': '\xe2\x9b\xb4',
	'field_hockey': '\xf0\x9f\x8f\x91',
	'fiji': '\xf0\x9f\x87\xab\xf0\x9f\x87\xaf',
	'file_cabinet': '\xf0\x9f\x97\x84',
	'file_folder': '\xf0\x9f\x93\x81',
	'film_projector': '\xf0\x9f\x93\xbd',
	'film_strip': '\xf0\x9f\x8e\x9e',
	'finland': '\xf0\x9f\x87\xab\xf0\x9f\x87\xae',
	'fire': '\xf0\x9f\x94\xa5',
	'fire_engine': '\xf0\x9f\x9a\x92',
	'fire_extinguisher': '\xf0\x9f\xa7\xaf',
	'firecracker': '\xf0\x9f\xa7\xa8',
	'firefighter': '\xf0\x9f\xa7\x91\xf0\x9f\x9a\x92',
	'fireworks': '\xf0\x9f\x8e\x86',
	'first_quarter_moon': '\xf0\x9f\x8c\x93',
	'first_quarter_moon_with_face': '\xf0\x9f\x8c\x9b',
	'fish': '\xf0\x9f\x90\x9f',
	'fish_cake': '\xf0\x9f\x8d\xa5',
	'fishing_pole_and_fish': '\xf0\x9f\x8e\xa3',
	'fist': '\xe2\x9c\x8a',
	'fist_left': '\xf0\x9f\xa4\x9b',
	'fist_oncoming': '\xf0\x9f\x91\x8a',
	'fist_raised': '\xe2\x9c\x8a',
	'fist_right': '\xf0\x9f\xa4\x9c',
	'five': '\x35\xe2\x83\xa3',
	'flags': '\xf0\x9f\x8e\x8f',
	'flamingo': '\xf0\x9f\xa6\xa9',
	'flashlight': '\xf0\x9f\x94\xa6',
	'flat_shoe': '\xf0\x9f\xa5\xbf',
	'flatbread': '\xf0\x9f\xab\x93',
	'fleur_de_lis': '\xe2\x9a\x9c',
	'flight_arrival': '\xf0\x9f\x9b\xac',
	'flight_departure': '\xf0\x9f\x9b\xab',
	'flipper': '\xf0\x9f\x90\xac',
	'floppy_disk': '\xf0\x9f\x92\xbe',
	'flower_playing_cards': '\xf0\x9f\x8e\xb4',
	'flushed': '\xf0\x9f\x98\xb3',
	'fly': '\xf0\x9f\xaa\xb0',
	'flying_disc': '\xf0\x9f\xa5\x8f',
	'flying_saucer': '\xf0\x9f\x9b\xb8',
	'fog': '\xf0\x9f\x8c\xab',
	'foggy': '\xf0\x9f\x8c\x81',
	'fondue': '\xf0\x9f\xab\x95',
	'foot': '\xf0\x9f\xa6\xb6',
	'football': '\xf0\x9f\x8f\x88',
	'footprints': '\xf0\x9f\x91\xa3',
	'fork_and_knife': '\xf0\x9f\x8d\xb4',
	'fortune_cookie': '\xf0\x9f\xa5\xa0',
	'fountain': '\xe2\x9b\xb2',
	'fountain_pen': '\xf0\x9f\x96\x8b',
	'four': '\x34\xe2\x83\xa3',
	'four_leaf_clover': '\xf0\x9f\x8d\x80',
	'fox_face': '\xf0\x9f\xa6\x8a',
	'fr': '\xf0\x9f\x87\xab\xf0\x9f\x87\xb7',
	'framed_picture': '\xf0\x9f\x96\xbc',
	'free': '\xf0\x9f\x86\x93',
	'french_guiana': '\xf0\x9f\x87\xac\xf0\x9f\x87\xab',
	'french_polynesia': '\xf0\x9f\x87\xb5\xf0\x9f\x87\xab',
	'french_southern_territories': '\xf0\x9f\x87\xb9\xf0\x9f\x87\xab',
	'fried_egg': '\xf0\x9f\x8d\xb3',
	'fried_shrimp': '\xf0\x9f\x8d\xa4',
	'fries': '\xf0\x9f\x8d\x9f',
	'frog': '\xf0\x9f\x90\xb8',
	'frowning': '\xf0\x9f\x98\xa6',
	'frowning_face': '\xe2\x98\xb9',
	'frowning_man': '\xf0\x9f\x99\x8d\xe2\x99\x82',
	'frowning_person': '\xf0\x9f\x99\x8d',
	'frowning_woman': '\xf0\x9f\x99\x8d\xe2\x99\x80',
	'fu': '\xf0\x9f\x96\x95',
	'fuelpump': '\xe2\x9b\xbd',
	'full_moon': '\xf0\x9f\x8c\x95',
	'full_moon_with_face': '\xf0\x9f\x8c\x9d',
	'funeral_urn': '\xe2\x9a\xb1',
	'gabon': '\xf0\x9f\x87\xac\xf0\x9f\x87\xa6',
	'gambia': '\xf0\x9f\x87\xac\xf0\x9f\x87\xb2',
	'game_die': '\xf0\x9f\x8e\xb2',
	'garlic': '\xf0\x9f\xa7\x84',
	'gb': '\xf0\x9f\x87\xac\xf0\x9f\x87\xa7',
	'gear': '\xe2\x9a\x99',
	'gem': '\xf0\x9f\x92\x8e',
	'gemini': '\xe2\x99\x8a',
	'genie': '\xf0\x9f\xa7\x9e',
	'genie_man': '\xf0\x9f\xa7\x9e\xe2\x99\x82',
	'genie_woman': '\xf0\x9f\xa7\x9e\xe2\x99\x80',
	'georgia': '\xf0\x9f\x87\xac\xf0\x9f\x87\xaa',
	'ghana': '\xf0\x9f\x87\xac\xf0\x9f\x87\xad',
	'ghost': '\xf0\x9f\x91\xbb',
	'gibraltar': '\xf0\x9f\x87\xac\xf0\x9f\x87\xae',
	'gift': '\xf0\x9f\x8e\x81',
	'gift_heart': '\xf0\x9f\x92\x9d',
	'giraffe': '\xf0\x9f\xa6\x92',
	'girl': '\xf0\x9f\x91\xa7',
	'globe_with_meridians': '\xf0\x9f\x8c\x90',
	'gloves': '\xf0\x9f\xa7\xa4',
	'goal_net': '\xf0\x9f\xa5\x85',
	'goat': '\xf0\x9f\x90\x90',
	'goggles': '\xf0\x9f\xa5\xbd',
	'golf': '\xe2\x9b\xb3',
	'golfing': '\xf0\x9f\x8f\x8c',
	'golfing_man': '\xf0\x9f\x8f\x8c\xe2\x99\x82',
	'golfing_woman': '\xf0\x9f\x8f\x8c\xe2\x99\x80',
	'gorilla': '\xf0\x9f\xa6\x8d',
	'grapes': '\xf0\x9f\x8d\x87',
	'greece': '\xf0\x9f\x87\xac\xf0\x9f\x87\xb7',
	'green_apple': '\xf0\x9f\x8d\x8f',
	'green_book': '\xf0\x9f\x93\x97',
	'green_circle': '\xf0\x9f\x9f\xa2',
	'green_heart': '\xf0\x9f\x92\x9a',
	'green_salad': '\xf0\x9f\xa5\x97',
	'green_square': '\xf0\x9f\x9f\xa9',
	'greenland': '\xf0\x9f\x87\xac\xf0\x9f\x87\xb1',
	'grenada': '\xf0\x9f\x87\xac\xf0\x9f\x87\xa9',
	'grey_exclamation': '\xe2\x9d\x95',
	'grey_question': '\xe2\x9d\x94',
	'grimacing': '\xf0\x9f\x98\xac',
	'grin': '\xf0\x9f\x98\x81',
	'grinning': '\xf0\x9f\x98\x80',
	'guadeloupe': '\xf0\x9f\x87\xac\xf0\x9f\x87\xb5',
	'guam': '\xf0\x9f\x87\xac\xf0\x9f\x87\xba',
	'guard': '\xf0\x9f\x92\x82',
	'guardsman': '\xf0\x9f\x92\x82\xe2\x99\x82',
	'guardswoman': '\xf0\x9f\x92\x82\xe2\x99\x80',
	'guatemala': '\xf0\x9f\x87\xac\xf0\x9f\x87\xb9',
	'guernsey': '\xf0\x9f\x87\xac\xf0\x9f\x87\xac',
	'guide_dog': '\xf0\x9f\xa6\xae',
	'guinea': '\xf0\x9f\x87\xac\xf0\x9f\x87\xb3',
	'guinea_bissau': '\xf0\x9f\x87\xac\xf0\x9f\x87\xbc',
	'guitar': '\xf0\x9f\x8e\xb8',
	'gun': '\xf0\x9f\x94\xab',
	'guyana': '\xf0\x9f\x87\xac\xf0\x9f\x87\xbe',
	'haircut': '\xf0\x9f\x92\x87',
	'haircut_man': '\xf0\x9f\x92\x87\xe2\x99\x82',
	'haircut_woman': '\xf0\x9f\x92\x87\xe2\x99\x80',
	'haiti': '\xf0\x9f\x87\xad\xf0\x9f\x87\xb9',
	'hamburger': '\xf0\x9f\x8d\x94',
	'hammer': '\xf0\x9f\x94\xa8',
	'hammer_and_pick': '\xe2\x9a\x92',
	'hammer_and_wrench': '\xf0\x9f\x9b\xa0',
	'hamster': '\xf0\x9f\x90\xb9',
	'hand': '\xe2\x9c\x8b',
	'hand_over_mouth': '\xf0\x9f\xa4\xad',
	'handbag': '\xf0\x9f\x91\x9c',
	'handball_person': '\xf0\x9f\xa4\xbe',
	'handshake': '\xf0\x9f\xa4\x9d',
	'hankey': '\xf0\x9f\x92\xa9',
	'hash': '\x23\xe2\x83\xa3',
	'hatched_chick': '\xf0\x9f\x90\xa5',
	'hatching_chick': '\xf0\x9f\x90\xa3',
	'headphones': '\xf0\x9f\x8e\xa7',
	'headstone': '\xf0\x9f\xaa\xa6',
	'health_worker': '\xf0\x9f\xa7\x91\xe2\x9a\x95',
	'hear_no_evil': '\xf0\x9f\x99\x89',
	'heard_mcdonald_islands': '\xf0\x9f\x87\xad\xf0\x9f\x87\xb2',
	'heart': '\xe2\x9d\xa4',
	'heart_decoration': '\xf0\x9f\x92\x9f',
	'heart_eyes': '\xf0\x9f\x98\x8d',
	'heart_eyes_cat': '\xf0\x9f\x98\xbb',
	'heart_on_fire': '\xe2\x9d\xa4\xf0\x9f\x94\xa5',
	'heartbeat': '\xf0\x9f\x92\x93',
	'heartpulse': '\xf0\x9f\x92\x97',
	'hearts': '\xe2\x99\xa5',
	'heavy_check_mark': '\xe2\x9c\x94',
	'heavy_division_sign': '\xe2\x9e\x97',
	'heavy_dollar_sign': '\xf0\x9f\x92\xb2',
	'heavy_exclamation_mark': '\xe2\x9d\x97',
	'heavy_heart_exclamation': '\xe2\x9d\xa3',
	'heavy_minus_sign': '\xe2\x9e\x96',
	'heavy_multiplication_x': '\xe2\x9c\x96',
	'heavy_plus_sign': '\xe2\x9e\x95',
	'hedgehog': '\xf0\x9f\xa6\x94',
	'helicopter': '\xf0\x9f\x9a\x81',
	'herb': '\xf0\x9f\x8c\xbf',
	'hibiscus': '\xf0\x9f\x8c\xba',
	'high_brightness': '\xf0\x9f\x94\x86',
	'high_heel': '\xf0\x9f\x91\xa0',
	'hiking_boot': '\xf0\x9f\xa5\xbe',
	'hindu_temple': '\xf0\x9f\x9b\x95',
	'hippopotamus': '\xf0\x9f\xa6\x9b',
	'hocho': '\xf0\x9f\x94\xaa',
	'hole': '\xf0\x9f\x95\xb3',
	'honduras': '\xf0\x9f\x87\xad\xf0\x9f\x87\xb3',
	'honey_pot': '\xf0\x9f\x8d\xaf',
	'honeybee': '\xf0\x9f\x90\x9d',
	'hong_kong': '\xf0\x9f\x87\xad\xf0\x9f\x87\xb0',
	'hook': '\xf0\x9f\xaa\x9d',
	'horse': '\xf0\x9f\x90\xb4',
	'horse_racing': '\xf0\x9f\x8f\x87',
	'hospital': '\xf0\x9f\x8f\xa5',
	'hot_face': '\xf0\x9f\xa5\xb5',
	'hot_pepper': '\xf0\x9f\x8c\xb6',
	'hotdog': '\xf0\x9f\x8c\xad',
	'hotel': '\xf0\x9f\x8f\xa8',
	'hotsprings': '\xe2\x99\xa8',
	'hourglass': '\xe2\x8c\x9b',
	'hourglass_flowing_sand': '\xe2\x8f\xb3',
	'house': '\xf0\x9f\x8f\xa0',
	'house_with_garden': '\xf0\x9f\x8f\xa1',
	'houses': '\xf0\x9f\x8f\x98',
	'hugs': '\xf0\x9f\xa4\x97',
	'hungary': '\xf0\x9f\x87\xad\xf0\x9f\x87\xba',
	'hushed': '\xf0\x9f\x98\xaf',
	'hut': '\xf0\x9f\x9b\x96',
	'ice_cream': '\xf0\x9f\x8d\xa8',
	'ice_cube': '\xf0\x9f\xa7\x8a',
	'ice_hockey': '\xf0\x9f\x8f\x92',
	'ice_skate': '\xe2\x9b\xb8',
	'icecream': '\xf0\x9f\x8d\xa6',
	'iceland': '\xf0\x9f\x87\xae\xf0\x9f\x87\xb8',
	'id': '\xf0\x9f\x86\x94',
	'ideograph_advantage': '\xf0\x9f\x89\x90',
	'imp': '\xf0\x9f\x91\xbf',
	'inbox_tray': '\xf0\x9f\x93\xa5',
	'incoming_envelope': '\xf0\x9f\x93\xa8',
	'india': '\xf0\x9f\x87\xae\xf0\x9f\x87\xb3',
	'indonesia': '\xf0\x9f\x87\xae\xf0\x9f\x87\xa9',
	'infinity': '\xe2\x99\xbe',
	'information_desk_person': '\xf0\x9f\x92\x81',
	'information_source': '\xe2\x84\xb9',
	'innocent': '\xf0\x9f\x98\x87',
	'interrobang': '\xe2\x81\x89',
	'iphone': '\xf0\x9f\x93\xb1',
	'iran': '\xf0\x9f\x87\xae\xf0\x9f\x87\xb7',
	'iraq': '\xf0\x9f\x87\xae\xf0\x9f\x87\xb6',
	'ireland': '\xf0\x9f\x87\xae\xf0\x9f\x87\xaa',
	'isle_of_man': '\xf0\x9f\x87\xae\xf0\x9f\x87\xb2',
	'israel': '\xf0\x9f\x87\xae\xf0\x9f\x87\xb1',
	'it': '\xf0\x9f\x87\xae\xf0\x9f\x87\xb9',
	'izakaya_lantern': '\xf0\x9f\x8f\xae',
	'jack_o_lantern': '\xf0\x9f\x8e\x83',
	'jamaica': '\xf0\x9f\x87\xaf\xf0\x9f\x87\xb2',
	'japan': '\xf0\x9f\x97\xbe',
	'japanese_castle': '\xf0\x9f\x8f\xaf',
	'japanese_goblin': '\xf0\x9f\x91\xba',
	'japanese_ogre': '\xf0\x9f\x91\xb9',
	'jeans': '\xf0\x9f\x91\x96',
	'jersey': '\xf0\x9f\x87\xaf\xf0\x9f\x87\xaa',
	'jigsaw': '\xf0\x9f\xa7\xa9',
	'jordan': '\xf0\x9f\x87\xaf\xf0\x9f\x87\xb4',
	'joy': '\xf0\x9f\x98\x82',
	'joy_cat': '\xf0\x9f\x98\xb9',
	'joystick': '\xf0\x9f\x95\xb9',
	'jp': '\xf0\x9f\x87\xaf\xf0\x9f\x87\xb5',
	'judge': '\xf0\x9f\xa7\x91\xe2\x9a\x96',
	'juggling_person': '\xf0\x9f\xa4\xb9',
	'kaaba': '\xf0\x9f\x95\x8b',
	'kangaroo': '\xf0\x9f\xa6\x98',
	'kazakhstan': '\xf0\x9f\x87\xb0\xf0\x9f\x87\xbf',
	'kenya': '\xf0\x9f\x87\xb0\xf0\x9f\x87\xaa',
	'key': '\xf0\x9f\x94\x91',
	'keyboard': '\xe2\x8c\xa8',
	'keycap_ten': '\xf0\x9f\x94\x9f',
	'kick_scooter': '\xf0\x9f\x9b\xb4',
	'kimono': '\xf0\x9f\x91\x98',
	'kiribati': '\xf0\x9f\x87\xb0\xf0\x9f\x87\xae',
	'kiss': '\xf0\x9f\x92\x8b',
	'kissing': '\xf0\x9f\x98\x97',
	'kissing_cat': '\xf0\x9f\x98\xbd',
	'kissing_closed_eyes': '\xf0\x9f\x98\x9a',
	'kissing_heart': '\xf0\x9f\x98\x98',
	'kissing_smiling_eyes': '\xf0\x9f\x98\x99',
	'kite': '\xf0\x9f\xaa\x81',
	'kiwi_fruit': '\xf0\x9f\xa5\x9d',
	'kneeling_man': '\xf0\x9f\xa7\x8e\xe2\x99\x82',
	'kneeling_person': '\xf0\x9f\xa7\x8e',
	'kneeling_woman': '\xf0\x9f\xa7\x8e\xe2\x99\x80',
	'knife': '\xf0\x9f\x94\xaa',
	'knot': '\xf0\x9f\xaa\xa2',
	'koala': '\xf0\x9f\x90\xa8',
	'koko': '\xf0\x9f\x88\x81',
	'kosovo': '\xf0\x9f\x87\xbd\xf0\x9f\x87\xb0',
	'kr': '\xf0\x9f\x87\xb0\xf0\x9f\x87\xb7',
	'kuwait': '\xf0\x9f\x87\xb0\xf0\x9f\x87\xbc',
	'kyrgyzstan': '\xf0\x9f\x87\xb0\xf0\x9f\x87\xac',
	'lab_coat': '\xf0\x9f\xa5\xbc',
	'label': '\xf0\x9f\x8f\xb7',
	'lacrosse': '\xf0\x9f\xa5\x8d',
	'ladder': '\xf0\x9f\xaa\x9c',
	'lady_beetle': '\xf0\x9f\x90\x9e',
	'lantern': '\xf0\x9f\x8f\xae',
	'laos': '\xf0\x9f\x87\xb1\xf0\x9f\x87\xa6',
	'large_blue_circle': '\xf0\x9f\x94\xb5',
	'large_blue_diamond': '\xf0\x9f\x94\xb7',
	'large_orange_diamond': '\xf0\x9f\x94\xb6',
	'last_quarter_moon': '\xf0\x9f\x8c\x97',
	'last_quarter_moon_with_face': '\xf0\x9f\x8c\x9c',
	'latin_cross': '\xe2\x9c\x9d',
	'latvia': '\xf0\x9f\x87\xb1\xf0\x9f\x87\xbb',
	'laughing': '\xf0\x9f\x98\x86',
	'leafy_green': '\xf0\x9f\xa5\xac',
	'leaves': '\xf0\x9f\x8d\x83',
	'lebanon': '\xf0\x9f\x87\xb1\xf0\x9f\x87\xa7',
	'ledger': '\xf0\x9f\x93\x92',
	'left_luggage': '\xf0\x9f\x9b\x85',
	'left_right_arrow': '\xe2\x86\x94',
	'left_speech_bubble': '\xf0\x9f\x97\xa8',
	'leftwards_arrow_with_hook': '\xe2\x86\xa9',
	'leg': '\xf0\x9f\xa6\xb5',
	'lemon': '\xf0\x9f\x8d\x8b',
	'leo': '\xe2\x99\x8c',
	'leopard': '\xf0\x9f\x90\x86',
	'lesotho': '\xf0\x9f\x87\xb1\xf0\x9f\x87\xb8',
	'level_slider': '\xf0\x9f\x8e\x9a',
	'liberia': '\xf0\x9f\x87\xb1\xf0\x9f\x87\xb7',
	'libra': '\xe2\x99\x8e',
	'libya': '\xf0\x9f\x87\xb1\xf0\x9f\x87\xbe',
	'liechtenstein': '\xf0\x9f\x87\xb1\xf0\x9f\x87\xae',
	'light_rail': '\xf0\x9f\x9a\x88',
	'link': '\xf0\x9f\x94\x97',
	'lion': '\xf0\x9f\xa6\x81',
	'lips': '\xf0\x9f\x91\x84',
	'lipstick': '\xf0\x9f\x92\x84',
	'lithuania': '\xf0\x9f\x87\xb1\xf0\x9f\x87\xb9',
	'lizard': '\xf0\x9f\xa6\x8e',
	'llama': '\xf0\x9f\xa6\x99',
	'lobster': '\xf0\x9f\xa6\x9e',
	'lock': '\xf0\x9f\x94\x92',
	'lock_with_ink_pen': '\xf0\x9f\x94\x8f',
	'lollipop': '\xf0\x9f\x8d\xad',
	'long_drum': '\xf0\x9f\xaa\x98',
	'loop': '\xe2\x9e\xbf',
	'lotion_bottle': '\xf0\x9f\xa7\xb4',
	'lotus_position': '\xf0\x9f\xa7\x98',
	'lotus_position_man': '\xf0\x9f\xa7\x98\xe2\x99\x82',
	'lotus_position_woman': '\xf0\x9f\xa7\x98\xe2\x99\x80',
	'loud_sound': '\xf0\x9f\x94\x8a',
	'loudspeaker': '\xf0\x9f\x93\xa2',
	'love_hotel': '\xf0\x9f\x8f\xa9',
	'love_letter': '\xf0\x9f\x92\x8c',
	'love_you_gesture': '\xf0\x9f\xa4\x9f',
	'low_brightness': '\xf0\x9f\x94\x85',
	'luggage': '\xf0\x9f\xa7\xb3',
	'lungs': '\xf0\x9f\xab\x81',
	'luxembourg': '\xf0\x9f\x87\xb1\xf0\x9f\x87\xba',
	'lying_face': '\xf0\x9f\xa4\xa5',
	'm': '\xe2\x93\x82',
	'macau': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xb4',
	'macedonia': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xb0',
	'madagascar': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xac',
	'mag': '\xf0\x9f\x94\x8d',
	'mag_right': '\xf0\x9f\x94\x8e',
	'mage': '\xf0\x9f\xa7\x99',
	'mage_man': '\xf0\x9f\xa7\x99\xe2\x99\x82',
	'mage_woman': '\xf0\x9f\xa7\x99\xe2\x99\x80',
	'magic_wand': '\xf0\x9f\xaa\x84',
	'magnet': '\xf0\x9f\xa7\xb2',
	'mahjong': '\xf0\x9f\x80\x84',
	'mailbox': '\xf0\x9f\x93\xab',
	'mailbox_closed': '\xf0\x9f\x93\xaa',
	'mailbox_with_mail': '\xf0\x9f\x93\xac',
	'mailbox_with_no_mail': '\xf0\x9f\x93\xad',
	'malawi': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xbc',
	'malaysia': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xbe',
	'maldives': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xbb',
	'male_detective': '\xf0\x9f\x95\xb5\xe2\x99\x82',
	'male_sign': '\xe2\x99\x82',
	'mali': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xb1',
	'malta': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xb9',
	'mammoth': '\xf0\x9f\xa6\xa3',
	'man': '\xf0\x9f\x91\xa8',
	'man_artist': '\xf0\x9f\x91\xa8\xf0\x9f\x8e\xa8',
	'man_astronaut': '\xf0\x9f\x91\xa8\xf0\x9f\x9a\x80',
	'man_beard': '\xf0\x9f\xa7\x94\xe2\x99\x82',
	'man_cartwheeling': '\xf0\x9f\xa4\xb8\xe2\x99\x82',
	'man_cook': '\xf0\x9f\x91\xa8\xf0\x9f\x8d\xb3',
	'man_dancing': '\xf0\x9f\x95\xba',
	'man_facepalming': '\xf0\x9f\xa4\xa6\xe2\x99\x82',
	'man_factory_worker': '\xf0\x9f\x91\xa8\xf0\x9f\x8f\xad',
	'man_farmer': '\xf0\x9f\x91\xa8\xf0\x9f\x8c\xbe',
	'man_feeding_baby': '\xf0\x9f\x91\xa8\xf0\x9f\x8d\xbc',
	'man_firefighter': '\xf0\x9f\x91\xa8\xf0\x9f\x9a\x92',
	'man_health_worker': '\xf0\x9f\x91\xa8\xe2\x9a\x95',
	'man_in_manual_wheelchair': '\xf0\x9f\x91\xa8\xf0\x9f\xa6\xbd',
	'man_in_motorized_wheelchair': '\xf0\x9f\x91\xa8\xf0\x9f\xa6\xbc',
	'man_in_tuxedo': '\xf0\x9f\xa4\xb5\xe2\x99\x82',
	'man_judge': '\xf0\x9f\x91\xa8\xe2\x9a\x96',
	'man_juggling': '\xf0\x9f\xa4\xb9\xe2\x99\x82',
	'man_mechanic': '\xf0\x9f\x91\xa8\xf0\x9f\x94\xa7',
	'man_office_worker': '\xf0\x9f\x91\xa8\xf0\x9f\x92\xbc',
	'man_pilot': '\xf0\x9f\x91\xa8\xe2\x9c\x88',
	'man_playing_handball': '\xf0\x9f\xa4\xbe\xe2\x99\x82',
	'man_playing_water_polo': '\xf0\x9f\xa4\xbd\xe2\x99\x82',
	'man_scientist': '\xf0\x9f\x91\xa8\xf0\x9f\x94\xac',
	'man_shrugging': '\xf0\x9f\xa4\xb7\xe2\x99\x82',
	'man_singer': '\xf0\x9f\x91\xa8\xf0\x9f\x8e\xa4',
	'man_student': '\xf0\x9f\x91\xa8\xf0\x9f\x8e\x93',
	'man_teacher': '\xf0\x9f\x91\xa8\xf0\x9f\x8f\xab',
	'man_technologist': '\xf0\x9f\x91\xa8\xf0\x9f\x92\xbb',
	'man_with_gua_pi_mao': '\xf0\x9f\x91\xb2',
	'man_with_probing_cane': '\xf0\x9f\x91\xa8\xf0\x9f\xa6\xaf',
	'man_with_turban': '\xf0\x9f\x91\xb3\xe2\x99\x82',
	'man_with_veil': '\xf0\x9f\x91\xb0\xe2\x99\x82',
	'mandarin': '\xf0\x9f\x8d\x8a',
	'mango': '\xf0\x9f\xa5\xad',
	'mans_shoe': '\xf0\x9f\x91\x9e',
	'mantelpiece_clock': '\xf0\x9f\x95\xb0',
	'manual_wheelchair': '\xf0\x9f\xa6\xbd',
	'maple_leaf': '\xf0\x9f\x8d\x81',
	'marshall_islands': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xad',
	'martial_arts_uniform': '\xf0\x9f\xa5\x8b',
	'martinique': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xb6',
	'mask': '\xf0\x9f\x98\xb7',
	'massage': '\xf0\x9f\x92\x86',
	'massage_man': '\xf0\x9f\x92\x86\xe2\x99\x82',
	'massage_woman': '\xf0\x9f\x92\x86\xe2\x99\x80',
	'mate': '\xf0\x9f\xa7\x89',
	'mauritania': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xb7',
	'mauritius': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xba',
	'mayotte': '\xf0\x9f\x87\xbe\xf0\x9f\x87\xb9',
	'meat_on_bone': '\xf0\x9f\x8d\x96',
	'mechanic': '\xf0\x9f\xa7\x91\xf0\x9f\x94\xa7',
	'mechanical_arm': '\xf0\x9f\xa6\xbe',
	'mechanical_leg': '\xf0\x9f\xa6\xbf',
	'medal_military': '\xf0\x9f\x8e\x96',
	'medal_sports': '\xf0\x9f\x8f\x85',
	'medical_symbol': '\xe2\x9a\x95',
	'mega': '\xf0\x9f\x93\xa3',
	'melon': '\xf0\x9f\x8d\x88',
	'memo': '\xf0\x9f\x93\x9d',
	'men_wrestling': '\xf0\x9f\xa4\xbc\xe2\x99\x82',
	'mending_heart': '\xe2\x9d\xa4\xf0\x9f\xa9\xb9',
	'menorah': '\xf0\x9f\x95\x8e',
	'mens': '\xf0\x9f\x9a\xb9',
	'mermaid': '\xf0\x9f\xa7\x9c\xe2\x99\x80',
	'merman': '\xf0\x9f\xa7\x9c\xe2\x99\x82',
	'merperson': '\xf0\x9f\xa7\x9c',
	'metal': '\xf0\x9f\xa4\x98',
	'metro': '\xf0\x9f\x9a\x87',
	'mexico': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xbd',
	'microbe': '\xf0\x9f\xa6\xa0',
	'micronesia': '\xf0\x9f\x87\xab\xf0\x9f\x87\xb2',
	'microphone': '\xf0\x9f\x8e\xa4',
	'microscope': '\xf0\x9f\x94\xac',
	'middle_finger': '\xf0\x9f\x96\x95',
	'military_helmet': '\xf0\x9f\xaa\x96',
	'milk_glass': '\xf0\x9f\xa5\x9b',
	'milky_way': '\xf0\x9f\x8c\x8c',
	'minibus': '\xf0\x9f\x9a\x90',
	'minidisc': '\xf0\x9f\x92\xbd',
	'mirror': '\xf0\x9f\xaa\x9e',
	'mobile_phone_off': '\xf0\x9f\x93\xb4',
	'moldova': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xa9',
	'monaco': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xa8',
	'money_mouth_face': '\xf0\x9f\xa4\x91',
	'money_with_wings': '\xf0\x9f\x92\xb8',
	'moneybag': '\xf0\x9f\x92\xb0',
	'mongolia': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xb3',
	'monkey': '\xf0\x9f\x90\x92',
	'monkey_face': '\xf0\x9f\x90\xb5',
	'monocle_face': '\xf0\x9f\xa7\x90',
	'monorail': '\xf0\x9f\x9a\x9d',
	'montenegro': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xaa',
	'montserrat': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xb8',
	'moon': '\xf0\x9f\x8c\x94',
	'moon_cake': '\xf0\x9f\xa5\xae',
	'morocco': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xa6',
	'mortar_board': '\xf0\x9f\x8e\x93',
	'mosque': '\xf0\x9f\x95\x8c',
	'mosquito': '\xf0\x9f\xa6\x9f',
	'motor_boat': '\xf0\x9f\x9b\xa5',
	'motor_scooter': '\xf0\x9f\x9b\xb5',
	'motorcycle': '\xf0\x9f\x8f\x8d',
	'motorized_wheelchair': '\xf0\x9f\xa6\xbc',
	'motorway': '\xf0\x9f\x9b\xa3',
	'mount_fuji': '\xf0\x9f\x97\xbb',
	'mountain': '\xe2\x9b\xb0',
	'mountain_bicyclist': '\xf0\x9f\x9a\xb5',
	'mountain_biking_man': '\xf0\x9f\x9a\xb5\xe2\x99\x82',
	'mountain_biking_woman': '\xf0\x9f\x9a\xb5\xe2\x99\x80',
	'mountain_cableway': '\xf0\x9f\x9a\xa0',
	'mountain_railway': '\xf0\x9f\x9a\x9e',
	'mountain_snow': '\xf0\x9f\x8f\x94',
	'mouse': '\xf0\x9f\x90\xad',
	'mouse2': '\xf0\x9f\x90\x81',
	'mouse_trap': '\xf0\x9f\xaa\xa4',
	'movie_camera': '\xf0\x9f\x8e\xa5',
	'moyai': '\xf0\x9f\x97\xbf',
	'mozambique': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xbf',
	'mrs_claus': '\xf0\x9f\xa4\xb6',
	'muscle': '\xf0\x9f\x92\xaa',
	'mushroom': '\xf0\x9f\x8d\x84',
	'musical_keyboard': '\xf0\x9f\x8e\xb9',
	'musical_note': '\xf0\x9f\x8e\xb5',
	'musical_score': '\xf0\x9f\x8e\xbc',
	'mute': '\xf0\x9f\x94\x87',
	'mx_claus': '\xf0\x9f\xa7\x91\xf0\x9f\x8e\x84',
	'myanmar': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xb2',
	'nail_care': '\xf0\x9f\x92\x85',
	'name_badge': '\xf0\x9f\x93\x9b',
	'namibia': '\xf0\x9f\x87\xb3\xf0\x9f\x87\xa6',
	'national_park': '\xf0\x9f\x8f\x9e',
	'nauru': '\xf0\x9f\x87\xb3\xf0\x9f\x87\xb7',
	'nauseated_face': '\xf0\x9f\xa4\xa2',
	'nazar_amulet': '\xf0\x9f\xa7\xbf',
	'necktie': '\xf0\x9f\x91\x94',
	'negative_squared_cross_mark': '\xe2\x9d\x8e',
	'nepal': '\xf0\x9f\x87\xb3\xf0\x9f\x87\xb5',
	'nerd_face': '\xf0\x9f\xa4\x93',
	'nesting_dolls': '\xf0\x9f\xaa\x86',
	'netherlands': '\xf0\x9f\x87\xb3\xf0\x9f\x87\xb1',
	'neutral_face': '\xf0\x9f\x98\x90',
	'new': '\xf0\x9f\x86\x95',
	'new_caledonia': '\xf0\x9f\x87\xb3\xf0\x9f\x87\xa8',
	'new_moon': '\xf0\x9f\x8c\x91',
	'new_moon_with_face': '\xf0\x9f\x8c\x9a',
	'new_zealand': '\xf0\x9f\x87\xb3\xf0\x9f\x87\xbf',
	'newspaper': '\xf0\x9f\x93\xb0',
	'newspaper_roll': '\xf0\x9f\x97\x9e',
	'next_track_button': '\xe2\x8f\xad',
	'ng': '\xf0\x9f\x86\x96',
	'ng_man': '\xf0\x9f\x99\x85\xe2\x99\x82',
	'ng_woman': '\xf0\x9f\x99\x85\xe2\x99\x80',
	'nicaragua': '\xf0\x9f\x87\xb3\xf0\x9f\x87\xae',
	'niger': '\xf0\x9f\x87\xb3\xf0\x9f\x87\xaa',
	'nigeria': '\xf0\x9f\x87\xb3\xf0\x9f\x87\xac',
	'night_with_stars': '\xf0\x9f\x8c\x83',
	'nine': '\x39\xe2\x83\xa3',
	'ninja': '\xf0\x9f\xa5\xb7',
	'niue': '\xf0\x9f\x87\xb3\xf0\x9f\x87\xba',
	'no_bell': '\xf0\x9f\x94\x95',
	'no_bicycles': '\xf0\x9f\x9a\xb3',
	'no_entry': '\xe2\x9b\x94',
	'no_entry_sign': '\xf0\x9f\x9a\xab',
	'no_good': '\xf0\x9f\x99\x85',
	'no_good_man': '\xf0\x9f\x99\x85\xe2\x99\x82',
	'no_good_woman': '\xf0\x9f\x99\x85\xe2\x99\x80',
	'no_mobile_phones': '\xf0\x9f\x93\xb5',
	'no_mouth': '\xf0\x9f\x98\xb6',
	'no_pedestrians': '\xf0\x9f\x9a\xb7',
	'no_smoking': '\xf0\x9f\x9a\xad',
	'non-potable_water': '\xf0\x9f\x9a\xb1',
	'norfolk_island': '\xf0\x9f\x87\xb3\xf0\x9f\x87\xab',
	'north_korea': '\xf0\x9f\x87\xb0\xf0\x9f\x87\xb5',
	'northern_mariana_islands': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xb5',
	'norway': '\xf0\x9f\x87\xb3\xf0\x9f\x87\xb4',
	'nose': '\xf0\x9f\x91\x83',
	'notebook': '\xf0\x9f\x93\x93',
	'notebook_with_decorative_cover': '\xf0\x9f\x93\x94',
	'notes': '\xf0\x9f\x8e\xb6',
	'nut_and_bolt': '\xf0\x9f\x94\xa9',
	'o': '\xe2\xad\x95',
	'o2': '\xf0\x9f\x85\xbe',
	'ocean': '\xf0\x9f\x8c\x8a',
	'octopus': '\xf0\x9f\x90\x99',
	'oden': '\xf0\x9f\x8d\xa2',
	'office': '\xf0\x9f\x8f\xa2',
	'office_worker': '\xf0\x9f\xa7\x91\xf0\x9f\x92\xbc',
	'oil_drum': '\xf0\x9f\x9b\xa2',
	'ok': '\xf0\x9f\x86\x97',
	'ok_hand': '\xf0\x9f\x91\x8c',
	'ok_man': '\xf0\x9f\x99\x86\xe2\x99\x82',
	'ok_person': '\xf0\x9f\x99\x86',
	'ok_woman': '\xf0\x9f\x99\x86\xe2\x99\x80',
	'old_key': '\xf0\x9f\x97\x9d',
	'older_adult': '\xf0\x9f\xa7\x93',
	'older_man': '\xf0\x9f\x91\xb4',
	'older_woman': '\xf0\x9f\x91\xb5',
	'olive': '\xf0\x9f\xab\x92',
	'om': '\xf0\x9f\x95\x89',
	'oman': '\xf0\x9f\x87\xb4\xf0\x9f\x87\xb2',
	'on': '\xf0\x9f\x94\x9b',
	'oncoming_automobile': '\xf0\x9f\x9a\x98',
	'oncoming_bus': '\xf0\x9f\x9a\x8d',
	'oncoming_police_car': '\xf0\x9f\x9a\x94',
	'oncoming_taxi': '\xf0\x9f\x9a\x96',
	'one': '\x31\xe2\x83\xa3',
	'one_piece_swimsuit': '\xf0\x9f\xa9\xb1',
	'onion': '\xf0\x9f\xa7\x85',
	'open_book': '\xf0\x9f\x93\x96',
	'open_file_folder': '\xf0\x9f\x93\x82',
	'open_hands': '\xf0\x9f\x91\x90',
	'open_mouth': '\xf0\x9f\x98\xae',
	'open_umbrella': '\xe2\x98\x82',
	'ophiuchus': '\xe2\x9b\x8e',
	'orange': '\xf0\x9f\x8d\x8a',
	'orange_book': '\xf0\x9f\x93\x99',
	'orange_circle': '\xf0\x9f\x9f\xa0',
	'orange_heart': '\xf0\x9f\xa7\xa1',
	'orange_square': '\xf0\x9f\x9f\xa7',
	'orangutan': '\xf0\x9f\xa6\xa7',
	'orthodox_cross': '\xe2\x98\xa6',
	'otter': '\xf0\x9f\xa6\xa6',
	'outbox_tray': '\xf0\x9f\x93\xa4',
	'owl': '\xf0\x9f\xa6\x89',
	'ox': '\xf0\x9f\x90\x82',
	'oyster': '\xf0\x9f\xa6\xaa',
	'package': '\xf0\x9f\x93\xa6',
	'page_facing_up': '\xf0\x9f\x93\x84',
	'page_with_curl': '\xf0\x9f\x93\x83',
	'pager': '\xf0\x9f\x93\x9f',
	'paintbrush': '\xf0\x9f\x96\x8c',
	'pakistan': '\xf0\x9f\x87\xb5\xf0\x9f\x87\xb0',
	'palau': '\xf0\x9f\x87\xb5\xf0\x9f\x87\xbc',
	'palestinian_territories': '\xf0\x9f\x87\xb5\xf0\x9f\x87\xb8',
	'palm_tree': '\xf0\x9f\x8c\xb4',
	'palms_up_together': '\xf0\x9f\xa4\xb2',
	'panama': '\xf0\x9f\x87\xb5\xf0\x9f\x87\xa6',
	'pancakes': '\xf0\x9f\xa5\x9e',
	'panda_face': '\xf0\x9f\x90\xbc',
	'paperclip': '\xf0\x9f\x93\x8e',
	'paperclips': '\xf0\x9f\x96\x87',
	'papua_new_guinea': '\xf0\x9f\x87\xb5\xf0\x9f\x87\xac',
	'parachute': '\xf0\x9f\xaa\x82',
	'paraguay': '\xf0\x9f\x87\xb5\xf0\x9f\x87\xbe',
	'parasol_on_ground': '\xe2\x9b\xb1',
	'parking': '\xf0\x9f\x85\xbf',
	'parrot': '\xf0\x9f\xa6\x9c',
	'part_alternation_mark': '\xe3\x80\xbd',
	'partly_sunny': '\xe2\x9b\x85',
	'partying_face': '\xf0\x9f\xa5\xb3',
	'passenger_ship': '\xf0\x9f\x9b\xb3',
	'passport_control': '\xf0\x9f\x9b\x82',
	'pause_button': '\xe2\x8f\xb8',
	'paw_prints': '\xf0\x9f\x90\xbe',
	'peace_symbol': '\xe2\x98\xae',
	'peach': '\xf0\x9f\x8d\x91',
	'peacock': '\xf0\x9f\xa6\x9a',
	'peanuts': '\xf0\x9f\xa5\x9c',
	'pear': '\xf0\x9f\x8d\x90',
	'pen': '\xf0\x9f\x96\x8a',
	'pencil': '\xf0\x9f\x93\x9d',
	'pencil2': '\xe2\x9c\x8f',
	'penguin': '\xf0\x9f\x90\xa7',
	'pensive': '\xf0\x9f\x98\x94',
	'people_holding_hands': '\xf0\x9f\xa7\x91\xf0\x9f\xa4\x9d\xf0\x9f\xa7\x91',
	'people_hugging': '\xf0\x9f\xab\x82',
	'performing_arts': '\xf0\x9f\x8e\xad',
	'persevere': '\xf0\x9f\x98\xa3',
	'person_bald': '\xf0\x9f\xa7\x91\xf0\x9f\xa6\xb2',
	'person_curly_hair': '\xf0\x9f\xa7\x91\xf0\x9f\xa6\xb1',
	'person_feeding_baby': '\xf0\x9f\xa7\x91\xf0\x9f\x8d\xbc',
	'person_fencing': '\xf0\x9f\xa4\xba',
	'person_in_manual_wheelchair': '\xf0\x9f\xa7\x91\xf0\x9f\xa6\xbd',
	'person_in_motorized_wheelchair': '\xf0\x9f\xa7\x91\xf0\x9f\xa6\xbc',
	'person_in_tuxedo': '\xf0\x9f\xa4\xb5',
	'person_red_hair': '\xf0\x9f\xa7\x91\xf0\x9f\xa6\xb0',
	'person_white_hair': '\xf0\x9f\xa7\x91\xf0\x9f\xa6\xb3',
	'person_with_probing_cane': '\xf0\x9f\xa7\x91\xf0\x9f\xa6\xaf',
	'person_with_turban': '\xf0\x9f\x91\xb3',
	'person_with_veil': '\xf0\x9f\x91\xb0',
	'peru': '\xf0\x9f\x87\xb5\xf0\x9f\x87\xaa',
	'petri_dish': '\xf0\x9f\xa7\xab',
	'philippines': '\xf0\x9f\x87\xb5\xf0\x9f\x87\xad',
	'phone': '\xe2\x98\x8e',
	'pick': '\xe2\x9b\x8f',
	'pickup_truck': '\xf0\x9f\x9b\xbb',
	'pie': '\xf0\x9f\xa5\xa7',
	'pig': '\xf0\x9f\x90\xb7',
	'pig2': '\xf0\x9f\x90\x96',
	'pig_nose': '\xf0\x9f\x90\xbd',
	'pill': '\xf0\x9f\x92\x8a',
	'pilot': '\xf0\x9f\xa7\x91\xe2\x9c\x88',
	'pinata': '\xf0\x9f\xaa\x85',
	'pinched_fingers': '\xf0\x9f\xa4\x8c',
	'pinching_hand': '\xf0\x9f\xa4\x8f',
	'pineapple': '\xf0\x9f\x8d\x8d',
	'ping_pong': '\xf0\x9f\x8f\x93',
	'pirate_flag': '\xf0\x9f\x8f\xb4\xe2\x98\xa0',
	'pisces': '\xe2\x99\x93',
	'pitcairn_islands': '\xf0\x9f\x87\xb5\xf0\x9f\x87\xb3',
	'pizza': '\xf0\x9f\x8d\x95',
	'placard': '\xf0\x9f\xaa\xa7',
	'place_of_worship': '\xf0\x9f\x9b\x90',
	'plate_with_cutlery': '\xf0\x9f\x8d\xbd',
	'play_or_pause_button': '\xe2\x8f\xaf',
	'pleading_face': '\xf0\x9f\xa5\xba',
	'plunger': '\xf0\x9f\xaa\xa0',
	'point_down': '\xf0\x9f\x91\x87',
	'point_left': '\xf0\x9f\x91\x88',
	'point_right': '\xf0\x9f\x91\x89',
	'point_up': '\xe2\x98\x9d',
	'point_up_2': '\xf0\x9f\x91\x86',
	'poland': '\xf0\x9f\x87\xb5\xf0\x9f\x87\xb1',
	'polar_bear': '\xf0\x9f\x90\xbb\xe2\x9d\x84',
	'police_car': '\xf0\x9f\x9a\x93',
	'police_officer': '\xf0\x9f\x91\xae',
	'policeman': '\xf0\x9f\x91\xae\xe2\x99\x82',
	'policewoman': '\xf0\x9f\x91\xae\xe2\x99\x80',
	'poodle': '\xf0\x9f\x90\xa9',
	'poop': '\xf0\x9f\x92\xa9',
	'popcorn': '\xf0\x9f\x8d\xbf',
	'portugal': '\xf0\x9f\x87\xb5\xf0\x9f\x87\xb9',
	'post_office': '\xf0\x9f\x8f\xa3',
	'postal_horn': '\xf0\x9f\x93\xaf',
	'postbox': '\xf0\x9f\x93\xae',
	'potable_water': '\xf0\x9f\x9a\xb0',
	'potato': '\xf0\x9f\xa5\x94',
	'potted_plant': '\xf0\x9f\xaa\xb4',
	'pouch': '\xf0\x9f\x91\x9d',
	'poultry_leg': '\xf0\x9f\x8d\x97',
	'pound': '\xf0\x9f\x92\xb7',
	'pout': '\xf0\x9f\x98\xa1',
	'pouting_cat': '\xf0\x9f\x98\xbe',
	'pouting_face': '\xf0\x9f\x99\x8e',
	'pouting_man': '\xf0\x9f\x99\x8e\xe2\x99\x82',
	'pouting_woman': '\xf0\x9f\x99\x8e\xe2\x99\x80',
	'pray': '\xf0\x9f\x99\x8f',
	'prayer_beads': '\xf0\x9f\x93\xbf',
	'pregnant_woman': '\xf0\x9f\xa4\xb0',
	'pretzel': '\xf0\x9f\xa5\xa8',
	'previous_track_button': '\xe2\x8f\xae',
	'prince': '\xf0\x9f\xa4\xb4',
	'princess': '\xf0\x9f\x91\xb8',
	'printer': '\xf0\x9f\x96\xa8',
	'probing_cane': '\xf0\x9f\xa6\xaf',
	'puerto_rico': '\xf0\x9f\x87\xb5\xf0\x9f\x87\xb7',
	'punch': '\xf0\x9f\x91\x8a',
	'purple_circle': '\xf0\x9f\x9f\xa3',
	'purple_heart': '\xf0\x9f\x92\x9c',
	'purple_square': '\xf0\x9f\x9f\xaa',
	'purse': '\xf0\x9f\x91\x9b',
	'pushpin': '\xf0\x9f\x93\x8c',
	'put_litter_in_its_place': '\xf0\x9f\x9a\xae',
	'qatar': '\xf0\x9f\x87\xb6\xf0\x9f\x87\xa6',
	'question': '\xe2\x9d\x93',
	'rabbit': '\xf0\x9f\x90\xb0',
	'rabbit2': '\xf0\x9f\x90\x87',
	'raccoon': '\xf0\x9f\xa6\x9d',
	'racehorse': '\xf0\x9f\x90\x8e',
	'racing_car': '\xf0\x9f\x8f\x8e',
	'radio': '\xf0\x9f\x93\xbb',
	'radio_button': '\xf0\x9f\x94\x98',
	'radioactive': '\xe2\x98\xa2',
	'rage': '\xf0\x9f\x98\xa1',
	'railway_car': '\xf0\x9f\x9a\x83',
	'railway_track': '\xf0\x9f\x9b\xa4',
	'rainbow': '\xf0\x9f\x8c\x88',
	'rainbow_flag': '\xf0\x9f\x8f\xb3\xf0\x9f\x8c\x88',
	'raised_back_of_hand': '\xf0\x9f\xa4\x9a',
	'raised_eyebrow': '\xf0\x9f\xa4\xa8',
	'raised_hand': '\xe2\x9c\x8b',
	'raised_hand_with_fingers_splayed': '\xf0\x9f\x96\x90',
	'raised_hands': '\xf0\x9f\x99\x8c',
	'raising_hand': '\xf0\x9f\x99\x8b',
	'raising_hand_man': '\xf0\x9f\x99\x8b\xe2\x99\x82',
	'raising_hand_woman': '\xf0\x9f\x99\x8b\xe2\x99\x80',
	'ram': '\xf0\x9f\x90\x8f',
	'ramen': '\xf0\x9f\x8d\x9c',
	'rat': '\xf0\x9f\x90\x80',
	'razor': '\xf0\x9f\xaa\x92',
	'receipt': '\xf0\x9f\xa7\xbe',
	'record_button': '\xe2\x8f\xba',
	'recycle': '\xe2\x99\xbb',
	'red_car': '\xf0\x9f\x9a\x97',
	'red_circle': '\xf0\x9f\x94\xb4',
	'red_envelope': '\xf0\x9f\xa7\xa7',
	'red_haired_man': '\xf0\x9f\x91\xa8\xf0\x9f\xa6\xb0',
	'red_haired_woman': '\xf0\x9f\x91\xa9\xf0\x9f\xa6\xb0',
	'red_square': '\xf0\x9f\x9f\xa5',
	'registered': '\xc2\xae',
	'relaxed': '\xe2\x98\xba',
	'relieved': '\xf0\x9f\x98\x8c',
	'reminder_ribbon': '\xf0\x9f\x8e\x97',
	'repeat': '\xf0\x9f\x94\x81',
	'repeat_one': '\xf0\x9f\x94\x82',
	'rescue_worker_helmet': '\xe2\x9b\x91',
	'restroom': '\xf0\x9f\x9a\xbb',
	'reunion': '\xf0\x9f\x87\xb7\xf0\x9f\x87\xaa',
	'revolving_hearts': '\xf0\x9f\x92\x9e',
	'rewind': '\xe2\x8f\xaa',
	'rhinoceros': '\xf0\x9f\xa6\x8f',
	'ribbon': '\xf0\x9f\x8e\x80',
	'rice': '\xf0\x9f\x8d\x9a',
	'rice_ball': '\xf0\x9f\x8d\x99',
	'rice_cracker': '\xf0\x9f\x8d\x98',
	'rice_scene': '\xf0\x9f\x8e\x91',
	'right_anger_bubble': '\xf0\x9f\x97\xaf',
	'ring': '\xf0\x9f\x92\x8d',
	'ringed_planet': '\xf0\x9f\xaa\x90',
	'robot': '\xf0\x9f\xa4\x96',
	'rock': '\xf0\x9f\xaa\xa8',
	'rocket': '\xf0\x9f\x9a\x80',
	'rofl': '\xf0\x9f\xa4\xa3',
	'roll_eyes': '\xf0\x9f\x99\x84',
	'roll_of_paper': '\xf0\x9f\xa7\xbb',
	'roller_coaster': '\xf0\x9f\x8e\xa2',
	'roller_skate': '\xf0\x9f\x9b\xbc',
	'romania': '\xf0\x9f\x87\xb7\xf0\x9f\x87\xb4',
	'rooster': '\xf0\x9f\x90\x93',
	'rose': '\xf0\x9f\x8c\xb9',
	'rosette': '\xf0\x9f\x8f\xb5',
	'rotating_light': '\xf0\x9f\x9a\xa8',
	'round_pushpin': '\xf0\x9f\x93\x8d',
	'rowboat': '\xf0\x9f\x9a\xa3',
	'rowing_man': '\xf0\x9f\x9a\xa3\xe2\x99\x82',
	'rowing_woman': '\xf0\x9f\x9a\xa3\xe2\x99\x80',
	'ru': '\xf0\x9f\x87\xb7\xf0\x9f\x87\xba',
	'rugby_football': '\xf0\x9f\x8f\x89',
	'runner': '\xf0\x9f\x8f\x83',
	'running': '\xf0\x9f\x8f\x83',
	'running_man': '\xf0\x9f\x8f\x83\xe2\x99\x82',
	'running_shirt_with_sash': '\xf0\x9f\x8e\xbd',
	'running_woman': '\xf0\x9f\x8f\x83\xe2\x99\x80',
	'rwanda': '\xf0\x9f\x87\xb7\xf0\x9f\x87\xbc',
	'sa': '\xf0\x9f\x88\x82',
	'safety_pin': '\xf0\x9f\xa7\xb7',
	'safety_vest': '\xf0\x9f\xa6\xba',
	'sagittarius': '\xe2\x99\x90',
	'sailboat': '\xe2\x9b\xb5',
	'sake': '\xf0\x9f\x8d\xb6',
	'salt': '\xf0\x9f\xa7\x82',
	'samoa': '\xf0\x9f\x87\xbc\xf0\x9f\x87\xb8',
	'san_marino': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xb2',
	'sandal': '\xf0\x9f\x91\xa1',
	'sandwich': '\xf0\x9f\xa5\xaa',
	'santa': '\xf0\x9f\x8e\x85',
	'sao_tome_principe': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xb9',
	'sari': '\xf0\x9f\xa5\xbb',
	'sassy_man': '\xf0\x9f\x92\x81\xe2\x99\x82',
	'sassy_woman': '\xf0\x9f\x92\x81\xe2\x99\x80',
	'satellite': '\xf0\x9f\x93\xa1',
	'satisfied': '\xf0\x9f\x98\x86',
	'saudi_arabia': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xa6',
	'sauna_man': '\xf0\x9f\xa7\x96\xe2\x99\x82',
	'sauna_person': '\xf0\x9f\xa7\x96',
	'sauna_woman': '\xf0\x9f\xa7\x96\xe2\x99\x80',
	'sauropod': '\xf0\x9f\xa6\x95',
	'saxophone': '\xf0\x9f\x8e\xb7',
	'scarf': '\xf0\x9f\xa7\xa3',
	'school': '\xf0\x9f\x8f\xab',
	'school_satchel': '\xf0\x9f\x8e\x92',
	'scientist': '\xf0\x9f\xa7\x91\xf0\x9f\x94\xac',
	'scissors': '\xe2\x9c\x82',
	'scorpion': '\xf0\x9f\xa6\x82',
	'scorpius': '\xe2\x99\x8f',
	'scotland': '\xf0\x9f\x8f\xb4\xf3\xa0\x81\xa7\xf3\xa0\x81\xa2\xf3\xa0\x81\xb3\xf3\xa0\x81\xa3\xf3\xa0\x81\xb4\xf3\xa0\x81\xbf',
	'scream': '\xf0\x9f\x98\xb1',
	'scream_cat': '\xf0\x9f\x99\x80',
	'screwdriver': '\xf0\x9f\xaa\x9b',
	'scroll': '\xf0\x9f\x93\x9c',
	'seal': '\xf0\x9f\xa6\xad',
	'seat': '\xf0\x9f\x92\xba',
	'secret': '\xe3\x8a\x99',
	'see_no_evil': '\xf0\x9f\x99\x88',
	'seedling': '\xf0\x9f\x8c\xb1',
	'selfie': '\xf0\x9f\xa4\xb3',
	'senegal': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xb3',
	'serbia': '\xf0\x9f\x87\xb7\xf0\x9f\x87\xb8',
	'service_dog': '\xf0\x9f\x90\x95\xf0\x9f\xa6\xba',
	'seven': '\x37\xe2\x83\xa3',
	'sewing_needle': '\xf0\x9f\xaa\xa1',
	'seychelles': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xa8',
	'shallow_pan_of_food': '\xf0\x9f\xa5\x98',
	'shamrock': '\xe2\x98\x98',
	'shark': '\xf0\x9f\xa6\x88',
	'shaved_ice': '\xf0\x9f\x8d\xa7',
	'sheep': '\xf0\x9f\x90\x91',
	'shell': '\xf0\x9f\x90\x9a',
	'shield': '\xf0\x9f\x9b\xa1',
	'shinto_shrine': '\xe2\x9b\xa9',
	'ship': '\xf0\x9f\x9a\xa2',
	'shirt': '\xf0\x9f\x91\x95',
	'shit': '\xf0\x9f\x92\xa9',
	'shoe': '\xf0\x9f\x91\x9e',
	'shopping': '\xf0\x9f\x9b\x8d',
	'shopping_cart': '\xf0\x9f\x9b\x92',
	'shorts': '\xf0\x9f\xa9\xb3',
	'shower': '\xf0\x9f\x9a\xbf',
	'shrimp': '\xf0\x9f\xa6\x90',
	'shrug': '\xf0\x9f\xa4\xb7',
	'shushing_face': '\xf0\x9f\xa4\xab',
	'sierra_leone': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xb1',
	'signal_strength': '\xf0\x9f\x93\xb6',
	'singapore': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xac',
	'singer': '\xf0\x9f\xa7\x91\xf0\x9f\x8e\xa4',
	'sint_maarten': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xbd',
	'six': '\x36\xe2\x83\xa3',
	'six_pointed_star': '\xf0\x9f\x94\xaf',
	'skateboard': '\xf0\x9f\x9b\xb9',
	'ski': '\xf0\x9f\x8e\xbf',
	'skier': '\xe2\x9b\xb7',
	'skull': '\xf0\x9f\x92\x80',
	'skull_and_crossbones': '\xe2\x98\xa0',
	'skunk': '\xf0\x9f\xa6\xa8',
	'sled': '\xf0\x9f\x9b\xb7',
	'sleeping': '\xf0\x9f\x98\xb4',
	'sleeping_bed': '\xf0\x9f\x9b\x8c',
	'sleepy': '\xf0\x9f\x98\xaa',
	'slightly_frowning_face': '\xf0\x9f\x99\x81',
	'slightly_smiling_face': '\xf0\x9f\x99\x82',
	'slot_machine': '\xf0\x9f\x8e\xb0',
	'sloth': '\xf0\x9f\xa6\xa5',
	'slovakia': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xb0',
	'slovenia': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xae',
	'small_airplane': '\xf0\x9f\x9b\xa9',
	'small_blue_diamond': '\xf0\x9f\x94\xb9',
	'small_orange_diamond': '\xf0\x9f\x94\xb8',
	'small_red_triangle': '\xf0\x9f\x94\xba',
	'small_red_triangle_down': '\xf0\x9f\x94\xbb',
	'smile': '\xf0\x9f\x98\x84',
	'smile_cat': '\xf0\x9f\x98\xb8',
	'smiley': '\xf0\x9f\x98\x83',
	'smiley_cat': '\xf0\x9f\x98\xba',
	'smiling_face_with_tear': '\xf0\x9f\xa5\xb2',
	'smiling_face_with_three_hearts': '\xf0\x9f\xa5\xb0',
	'smiling_imp': '\xf0\x9f\x98\x88',
	'smirk': '\xf0\x9f\x98\x8f',
	'smirk_cat': '\xf0\x9f\x98\xbc',
	'smoking': '\xf0\x9f\x9a\xac',
	'snail': '\xf0\x9f\x90\x8c',
	'snake': '\xf0\x9f\x90\x8d',
	'sneezing_face': '\xf0\x9f\xa4\xa7',
	'snowboarder': '\xf0\x9f\x8f\x82',
	'snowflake': '\xe2\x9d\x84',
	'snowman': '\xe2\x9b\x84',
	'snowman_with_snow': '\xe2\x98\x83',
	'soap': '\xf0\x9f\xa7\xbc',
	'sob': '\xf0\x9f\x98\xad',
	'soccer': '\xe2\x9a\xbd',
	'socks': '\xf0\x9f\xa7\xa6',
	'softball': '\xf0\x9f\xa5\x8e',
	'solomon_islands': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xa7',
	'somalia': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xb4',
	'soon': '\xf0\x9f\x94\x9c',
	'sos': '\xf0\x9f\x86\x98',
	'sound': '\xf0\x9f\x94\x89',
	'south_africa': '\xf0\x9f\x87\xbf\xf0\x9f\x87\xa6',
	'south_georgia_south_sandwich_islands': '\xf0\x9f\x87\xac\xf0\x9f\x87\xb8',
	'south_sudan': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xb8',
	'space_invader': '\xf0\x9f\x91\xbe',
	'spades': '\xe2\x99\xa0',
	'spaghetti': '\xf0\x9f\x8d\x9d',
	'sparkle': '\xe2\x9d\x87',
	'sparkler': '\xf0\x9f\x8e\x87',
	'sparkles': '\xe2\x9c\xa8',
	'sparkling_heart': '\xf0\x9f\x92\x96',
	'speak_no_evil': '\xf0\x9f\x99\x8a',
	'speaker': '\xf0\x9f\x94\x88',
	'speaking_head': '\xf0\x9f\x97\xa3',
	'speech_balloon': '\xf0\x9f\x92\xac',
	'speedboat': '\xf0\x9f\x9a\xa4',
	'spider': '\xf0\x9f\x95\xb7',
	'spider_web': '\xf0\x9f\x95\xb8',
	'spiral_calendar': '\xf0\x9f\x97\x93',
	'spiral_notepad': '\xf0\x9f\x97\x92',
	'sponge': '\xf0\x9f\xa7\xbd',
	'spoon': '\xf0\x9f\xa5\x84',
	'squid': '\xf0\x9f\xa6\x91',
	'sri_lanka': '\xf0\x9f\x87\xb1\xf0\x9f\x87\xb0',
	'st_barthelemy': '\xf0\x9f\x87\xa7\xf0\x9f\x87\xb1',
	'st_helena': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xad',
	'st_kitts_nevis': '\xf0\x9f\x87\xb0\xf0\x9f\x87\xb3',
	'st_lucia': '\xf0\x9f\x87\xb1\xf0\x9f\x87\xa8',
	'st_martin': '\xf0\x9f\x87\xb2\xf0\x9f\x87\xab',
	'st_pierre_miquelon': '\xf0\x9f\x87\xb5\xf0\x9f\x87\xb2',
	'st_vincent_grenadines': '\xf0\x9f\x87\xbb\xf0\x9f\x87\xa8',
	'stadium': '\xf0\x9f\x8f\x9f',
	'standing_man': '\xf0\x9f\xa7\x8d\xe2\x99\x82',
	'standing_person': '\xf0\x9f\xa7\x8d',
	'standing_woman': '\xf0\x9f\xa7\x8d\xe2\x99\x80',
	'star': '\xe2\xad\x90',
	'star2': '\xf0\x9f\x8c\x9f',
	'star_and_crescent': '\xe2\x98\xaa',
	'star_of_david': '\xe2\x9c\xa1',
	'star_struck': '\xf0\x9f\xa4\xa9',
	'stars': '\xf0\x9f\x8c\xa0',
	'station': '\xf0\x9f\x9a\x89',
	'statue_of_liberty': '\xf0\x9f\x97\xbd',
	'steam_locomotive': '\xf0\x9f\x9a\x82',
	'stethoscope': '\xf0\x9f\xa9\xba',
	'stew': '\xf0\x9f\x8d\xb2',
	'stop_button': '\xe2\x8f\xb9',
	'stop_sign': '\xf0\x9f\x9b\x91',
	'stopwatch': '\xe2\x8f\xb1',
	'straight_ruler': '\xf0\x9f\x93\x8f',
	'strawberry': '\xf0\x9f\x8d\x93',
	'stuck_out_tongue': '\xf0\x9f\x98\x9b',
	'stuck_out_tongue_closed_eyes': '\xf0\x9f\x98\x9d',
	'stuck_out_tongue_winking_eye': '\xf0\x9f\x98\x9c',
	'student': '\xf0\x9f\xa7\x91\xf0\x9f\x8e\x93',
	'studio_microphone': '\xf0\x9f\x8e\x99',
	'stuffed_flatbread': '\xf0\x9f\xa5\x99',
	'sudan': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xa9',
	'sun_behind_large_cloud': '\xf0\x9f\x8c\xa5',
	'sun_behind_rain_cloud': '\xf0\x9f\x8c\xa6',
	'sun_behind_small_cloud': '\xf0\x9f\x8c\xa4',
	'sun_with_face': '\xf0\x9f\x8c\x9e',
	'sunflower': '\xf0\x9f\x8c\xbb',
	'sunglasses': '\xf0\x9f\x98\x8e',
	'sunny': '\xe2\x98\x80',
	'sunrise': '\xf0\x9f\x8c\x85',
	'sunrise_over_mountains': '\xf0\x9f\x8c\x84',
	'superhero': '\xf0\x9f\xa6\xb8',
	'superhero_man': '\xf0\x9f\xa6\xb8\xe2\x99\x82',
	'superhero_woman': '\xf0\x9f\xa6\xb8\xe2\x99\x80',
	'supervillain': '\xf0\x9f\xa6\xb9',
	'supervillain_man': '\xf0\x9f\xa6\xb9\xe2\x99\x82',
	'supervillain_woman': '\xf0\x9f\xa6\xb9\xe2\x99\x80',
	'surfer': '\xf0\x9f\x8f\x84',
	'surfing_man': '\xf0\x9f\x8f\x84\xe2\x99\x82',
	'surfing_woman': '\xf0\x9f\x8f\x84\xe2\x99\x80',
	'suriname': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xb7',
	'sushi': '\xf0\x9f\x8d\xa3',
	'suspension_railway': '\xf0\x9f\x9a\x9f',
	'svalbard_jan_mayen': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xaf',
	'swan': '\xf0\x9f\xa6\xa2',
	'swaziland': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xbf',
	'sweat': '\xf0\x9f\x98\x93',
	'sweat_drops': '\xf0\x9f\x92\xa6',
	'sweat_smile': '\xf0\x9f\x98\x85',
	'sweden': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xaa',
	'sweet_potato': '\xf0\x9f\x8d\xa0',
	'swim_brief': '\xf0\x9f\xa9\xb2',
	'swimmer': '\xf0\x9f\x8f\x8a',
	'swimming_man': '\xf0\x9f\x8f\x8a\xe2\x99\x82',
	'swimming_woman': '\xf0\x9f\x8f\x8a\xe2\x99\x80',
	'switzerland': '\xf0\x9f\x87\xa8\xf0\x9f\x87\xad',
	'symbols': '\xf0\x9f\x94\xa3',
	'synagogue': '\xf0\x9f\x95\x8d',
	'syria': '\xf0\x9f\x87\xb8\xf0\x9f\x87\xbe',
	'syringe': '\xf0\x9f\x92\x89',
	't-rex': '\xf0\x9f\xa6\x96',
	'taco': '\xf0\x9f\x8c\xae',
	'tada': '\xf0\x9f\x8e\x89',
	'taiwan': '\xf0\x9f\x87\xb9\xf0\x9f\x87\xbc',
	'tajikistan': '\xf0\x9f\x87\xb9\xf0\x9f\x87\xaf',
	'takeout_box': '\xf0\x9f\xa5\xa1',
	'tamale': '\xf0\x9f\xab\x94',
	'tanabata_tree': '\xf0\x9f\x8e\x8b',
	'tangerine': '\xf0\x9f\x8d\x8a',
	'tanzania': '\xf0\x9f\x87\xb9\xf0\x9f\x87\xbf',
	'taurus': '\xe2\x99\x89',
	'taxi': '\xf0\x9f\x9a\x95',
	'tea': '\xf0\x9f\x8d\xb5',
	'teacher': '\xf0\x9f\xa7\x91\xf0\x9f\x8f\xab',
	'teapot': '\xf0\x9f\xab\x96',
	'technologist': '\xf0\x9f\xa7\x91\xf0\x9f\x92\xbb',
	'teddy_bear': '\xf0\x9f\xa7\xb8',
	'telephone': '\xe2\x98\x8e',
	'telephone_receiver': '\xf0\x9f\x93\x9e',
	'telescope': '\xf0\x9f\x94\xad',
	'tennis': '\xf0\x9f\x8e\xbe',
	'tent': '\xe2\x9b\xba',
	'test_tube': '\xf0\x9f\xa7\xaa',
	'thailand': '\xf0\x9f\x87\xb9\xf0\x9f\x87\xad',
	'thermometer': '\xf0\x9f\x8c\xa1',
	'thinking': '\xf0\x9f\xa4\x94',
	'thong_sandal': '\xf0\x9f\xa9\xb4',
	'thought_balloon': '\xf0\x9f\x92\xad',
	'thread': '\xf0\x9f\xa7\xb5',
	'three': '\x33\xe2\x83\xa3',
	'thumbsdown': '\xf0\x9f\x91\x8e',
	'thumbsup': '\xf0\x9f\x91\x8d',
	'ticket': '\xf0\x9f\x8e\xab',
	'tickets': '\xf0\x9f\x8e\x9f',
	'tiger': '\xf0\x9f\x90\xaf',
	'tiger2': '\xf0\x9f\x90\x85',
	'timer_clock': '\xe2\x8f\xb2',
	'timor_leste': '\xf0\x9f\x87\xb9\xf0\x9f\x87\xb1',
	'tipping_hand_man': '\xf0\x9f\x92\x81\xe2\x99\x82',
	'tipping_hand_person': '\xf0\x9f\x92\x81',
	'tipping_hand_woman': '\xf0\x9f\x92\x81\xe2\x99\x80',
	'tired_face': '\xf0\x9f\x98\xab',
	'tm': '\xe2\x84\xa2',
	'togo': '\xf0\x9f\x87\xb9\xf0\x9f\x87\xac',
	'toilet': '\xf0\x9f\x9a\xbd',
	'tokelau': '\xf0\x9f\x87\xb9\xf0\x9f\x87\xb0',
	'tokyo_tower': '\xf0\x9f\x97\xbc',
	'tomato': '\xf0\x9f\x8d\x85',
	'tonga': '\xf0\x9f\x87\xb9\xf0\x9f\x87\xb4',
	'tongue': '\xf0\x9f\x91\x85',
	'toolbox': '\xf0\x9f\xa7\xb0',
	'tooth': '\xf0\x9f\xa6\xb7',
	'toothbrush': '\xf0\x9f\xaa\xa5',
	'top': '\xf0\x9f\x94\x9d',
	'tophat': '\xf0\x9f\x8e\xa9',
	'tornado': '\xf0\x9f\x8c\xaa',
	'tr': '\xf0\x9f\x87\xb9\xf0\x9f\x87\xb7',
	'trackball': '\xf0\x9f\x96\xb2',
	'tractor': '\xf0\x9f\x9a\x9c',
	'traffic_light': '\xf0\x9f\x9a\xa5',
	'train': '\xf0\x9f\x9a\x8b',
	'train2': '\xf0\x9f\x9a\x86',
	'tram': '\xf0\x9f\x9a\x8a',
	'transgender_flag': '\xf0\x9f\x8f\xb3\xe2\x9a\xa7',
	'transgender_symbol': '\xe2\x9a\xa7',
	'triangular_flag_on_post': '\xf0\x9f\x9a\xa9',
	'triangular_ruler': '\xf0\x9f\x93\x90',
	'trident': '\xf0\x9f\x94\xb1',
	'trinidad_tobago': '\xf0\x9f\x87\xb9\xf0\x9f\x87\xb9',
	'tristan_da_cunha': '\xf0\x9f\x87\xb9\xf0\x9f\x87\xa6',
	'triumph': '\xf0\x9f\x98\xa4',
	'trolleybus': '\xf0\x9f\x9a\x8e',
	'trophy': '\xf0\x9f\x8f\x86',
	'tropical_drink': '\xf0\x9f\x8d\xb9',
	'tropical_fish': '\xf0\x9f\x90\xa0',
	'truck': '\xf0\x9f\x9a\x9a',
	'trumpet': '\xf0\x9f\x8e\xba',
	'tshirt': '\xf0\x9f\x91\x95',
	'tulip': '\xf0\x9f\x8c\xb7',
	'tumbler_glass': '\xf0\x9f\xa5\x83',
	'tunisia': '\xf0\x9f\x87\xb9\xf0\x9f\x87\xb3',
	'turkey': '\xf0\x9f\xa6\x83',
	'turkmenistan': '\xf0\x9f\x87\xb9\xf0\x9f\x87\xb2',
	'turks_caicos_islands': '\xf0\x9f\x87\xb9\xf0\x9f\x87\xa8',
	'turtle': '\xf0\x9f\x90\xa2',
	'tuvalu': '\xf0\x9f\x87\xb9\xf0\x9f\x87\xbb',
	'tv': '\xf0\x9f\x93\xba',
	'twisted_rightwards_arrows': '\xf0\x9f\x94\x80',
	'two': '\x32\xe2\x83\xa3',
	'two_hearts': '\xf0\x9f\x92\x95',
	'two_men_holding_hands': '\xf0\x9f\x91\xac',
	'two_women_holding_hands': '\xf0\x9f\x91\xad',
	'u5272': '\xf0\x9f\x88\xb9',
	'u5408': '\xf0\x9f\x88\xb4',
	'u55b6': '\xf0\x9f\x88\xba',
	'u6307': '\xf0\x9f\x88\xaf',
	'u6708': '\xf0\x9f\x88\xb7',
	'u6709': '\xf0\x9f\x88\xb6',
	'u6e80': '\xf0\x9f\x88\xb5',
	'u7121': '\xf0\x9f\x88\x9a',
	'u7533': '\xf0\x9f\x88\xb8',
	'u7981': '\xf0\x9f\x88\xb2',
	'u7a7a': '\xf0\x9f\x88\xb3',
	'uganda': '\xf0\x9f\x87\xba\xf0\x9f\x87\xac',
	'uk': '\xf0\x9f\x87\xac\xf0\x9f\x87\xa7',
	'ukraine': '\xf0\x9f\x87\xba\xf0\x9f\x87\xa6',
	'umbrella': '\xe2\x98\x94',
	'unamused': '\xf0\x9f\x98\x92',
	'underage': '\xf0\x9f\x94\x9e',
	'unicorn': '\xf0\x9f\xa6\x84',
	'united_arab_emirates': '\xf0\x9f\x87\xa6\xf0\x9f\x87\xaa',
	'united_nations': '\xf0\x9f\x87\xba\xf0\x9f\x87\xb3',
	'unlock': '\xf0\x9f\x94\x93',
	'up': '\xf0\x9f\x86\x99',
	'upside_down_face': '\xf0\x9f\x99\x83',
	'uruguay': '\xf0\x9f\x87\xba\xf0\x9f\x87\xbe',
	'us': '\xf0\x9f\x87\xba\xf0\x9f\x87\xb8',
	'us_outlying_islands': '\xf0\x9f\x87\xba\xf0\x9f\x87\xb2',
	'us_virgin_islands': '\xf0\x9f\x87\xbb\xf0\x9f\x87\xae',
	'uzbekistan': '\xf0\x9f\x87\xba\xf0\x9f\x87\xbf',
	'v': '\xe2\x9c\x8c',
	'vampire': '\xf0\x9f\xa7\x9b',
	'vampire_man': '\xf0\x9f\xa7\x9b\xe2\x99\x82',
	'vampire_woman': '\xf0\x9f\xa7\x9b\xe2\x99\x80',
	'vanuatu': '\xf0\x9f\x87\xbb\xf0\x9f\x87\xba',
	'vatican_city': '\xf0\x9f\x87\xbb\xf0\x9f\x87\xa6',
	'venezuela': '\xf0\x9f\x87\xbb\xf0\x9f\x87\xaa',
	'vertical_traffic_light': '\xf0\x9f\x9a\xa6',
	'vhs': '\xf0\x9f\x93\xbc',
	'vibration_mode': '\xf0\x9f\x93\xb3',
	'video_camera': '\xf0\x9f\x93\xb9',
	'video_game': '\xf0\x9f\x8e\xae',
	'vietnam': '\xf0\x9f\x87\xbb\xf0\x9f\x87\xb3',
	'violin': '\xf0\x9f\x8e\xbb',
	'virgo': '\xe2\x99\x8d',
	'volcano': '\xf0\x9f\x8c\x8b',
	'volleyball': '\xf0\x9f\x8f\x90',
	'vomiting_face': '\xf0\x9f\xa4\xae',
	'vs': '\xf0\x9f\x86\x9a',
	'vulcan_salute': '\xf0\x9f\x96\x96',
	'waffle': '\xf0\x9f\xa7\x87',
	'wales': '\xf0\x9f\x8f\xb4\xf3\xa0\x81\xa7\xf3\xa0\x81\xa2\xf3\xa0\x81\xb7\xf3\xa0\x81\xac\xf3\xa0\x81\xb3\xf3\xa0\x81\xbf',
	'walking': '\xf0\x9f\x9a\xb6',
	'walking_man': '\xf0\x9f\x9a\xb6\xe2\x99\x82',
	'walking_woman': '\xf0\x9f\x9a\xb6\xe2\x99\x80',
	'wallis_futuna': '\xf0\x9f\x87\xbc\xf0\x9f\x87\xab',
	'waning_crescent_moon': '\xf0\x9f\x8c\x98',
	'waning_gibbous_moon': '\xf0\x9f\x8c\x96',
	'warning': '\xe2\x9a\xa0',
	'wastebasket': '\xf0\x9f\x97\x91',
	'watch': '\xe2\x8c\x9a',
	'water_buffalo': '\xf0\x9f\x90\x83',
	'water_polo': '\xf0\x9f\xa4\xbd',
	'watermelon': '\xf0\x9f\x8d\x89',
	'wave': '\xf0\x9f\x91\x8b',
	'wavy_dash': '\xe3\x80\xb0',
	'waxing_crescent_moon': '\xf0\x9f\x8c\x92',
	'waxing_gibbous_moon': '\xf0\x9f\x8c\x94',
	'wc': '\xf0\x9f\x9a\xbe',
	'weary': '\xf0\x9f\x98\xa9',
	'wedding': '\xf0\x9f\x92\x92',
	'weight_lifting': '\xf0\x9f\x8f\x8b',
	'weight_lifting_man': '\xf0\x9f\x8f\x8b\xe2\x99\x82',
	'weight_lifting_woman': '\xf0\x9f\x8f\x8b\xe2\x99\x80',
	'western_sahara': '\xf0\x9f\x87\xaa\xf0\x9f\x87\xad',
	'whale': '\xf0\x9f\x90\xb3',
	'whale2': '\xf0\x9f\x90\x8b',
	'wheel_of_dharma': '\xe2\x98\xb8',
	'wheelchair': '\xe2\x99\xbf',
	'white_check_mark': '\xe2\x9c\x85',
	'white_circle': '\xe2\x9a\xaa',
	'white_flag': '\xf0\x9f\x8f\xb3',
	'white_flower': '\xf0\x9f\x92\xae',
	'white_haired_man': '\xf0\x9f\x91\xa8\xf0\x9f\xa6\xb3',
	'white_haired_woman': '\xf0\x9f\x91\xa9\xf0\x9f\xa6\xb3',
	'white_heart': '\xf0\x9f\xa4\x8d',
	'white_large_square': '\xe2\xac\x9c',
	'white_medium_small_square': '\xe2\x97\xbd',
	'white_medium_square': '\xe2\x97\xbb',
	'white_small_square': '\xe2\x96\xab',
	'white_square_button': '\xf0\x9f\x94\xb3',
	'wilted_flower': '\xf0\x9f\xa5\x80',
	'wind_chime': '\xf0\x9f\x8e\x90',
	'wind_face': '\xf0\x9f\x8c\xac',
	'window': '\xf0\x9f\xaa\x9f',
	'wine_glass': '\xf0\x9f\x8d\xb7',
	'wink': '\xf0\x9f\x98\x89',
	'wolf': '\xf0\x9f\x90\xba',
	'woman': '\xf0\x9f\x91\xa9',
	'woman_artist': '\xf0\x9f\x91\xa9\xf0\x9f\x8e\xa8',
	'woman_astronaut': '\xf0\x9f\x91\xa9\xf0\x9f\x9a\x80',
	'woman_beard': '\xf0\x9f\xa7\x94\xe2\x99\x80',
	'woman_cartwheeling': '\xf0\x9f\xa4\xb8\xe2\x99\x80',
	'woman_cook': '\xf0\x9f\x91\xa9\xf0\x9f\x8d\xb3',
	'woman_dancing': '\xf0\x9f\x92\x83',
	'woman_facepalming': '\xf0\x9f\xa4\xa6\xe2\x99\x80',
	'woman_factory_worker': '\xf0\x9f\x91\xa9\xf0\x9f\x8f\xad',
	'woman_farmer': '\xf0\x9f\x91\xa9\xf0\x9f\x8c\xbe',
	'woman_feeding_baby': '\xf0\x9f\x91\xa9\xf0\x9f\x8d\xbc',
	'woman_firefighter': '\xf0\x9f\x91\xa9\xf0\x9f\x9a\x92',
	'woman_health_worker': '\xf0\x9f\x91\xa9\xe2\x9a\x95',
	'woman_in_manual_wheelchair': '\xf0\x9f\x91\xa9\xf0\x9f\xa6\xbd',
	'woman_in_motorized_wheelchair': '\xf0\x9f\x91\xa9\xf0\x9f\xa6\xbc',
	'woman_in_tuxedo': '\xf0\x9f\xa4\xb5\xe2\x99\x80',
	'woman_judge': '\xf0\x9f\x91\xa9\xe2\x9a\x96',
	'woman_juggling': '\xf0\x9f\xa4\xb9\xe2\x99\x80',
	'woman_mechanic': '\xf0\x9f\x91\xa9\xf0\x9f\x94\xa7',
	'woman_office_worker': '\xf0\x9f\x91\xa9\xf0\x9f\x92\xbc',
	'woman_pilot': '\xf0\x9f\x91\xa9\xe2\x9c\x88',
	'woman_playing_handball': '\xf0\x9f\xa4\xbe\xe2\x99\x80',
	'woman_playing_water_polo': '\xf0\x9f\xa4\xbd\xe2\x99\x80',
	'woman_scientist': '\xf0\x9f\x91\xa9\xf0\x9f\x94\xac',
	'woman_shrugging': '\xf0\x9f\xa4\xb7\xe2\x99\x80',
	'woman_singer': '\xf0\x9f\x91\xa9\xf0\x9f\x8e\xa4',
	'woman_student': '\xf0\x9f\x91\xa9\xf0\x9f\x8e\x93',
	'woman_teacher': '\xf0\x9f\x91\xa9\xf0\x9f\x8f\xab',
	'woman_technologist': '\xf0\x9f\x91\xa9\xf0\x9f\x92\xbb',
	'woman_with_headscarf': '\xf0\x9f\xa7\x95',
	'woman_with_probing_cane': '\xf0\x9f\x91\xa9\xf0\x9f\xa6\xaf',
	'woman_with_turban': '\xf0\x9f\x91\xb3\xe2\x99\x80',
	'woman_with_veil': '\xf0\x9f\x91\xb0\xe2\x99\x80',
	'womans_clothes': '\xf0\x9f\x91\x9a',
	'womans_hat': '\xf0\x9f\x91\x92',
	'women_wrestling': '\xf0\x9f\xa4\xbc\xe2\x99\x80',
	'womens': '\xf0\x9f\x9a\xba',
	'wood': '\xf0\x9f\xaa\xb5',
	'woozy_face': '\xf0\x9f\xa5\xb4',
	'world_map': '\xf0\x9f\x97\xba',
	'worm': '\xf0\x9f\xaa\xb1',
	'worried': '\xf0\x9f\x98\x9f',
	'wrench': '\xf0\x9f\x94\xa7',
	'wrestling': '\xf0\x9f\xa4\xbc',
	'writing_hand': '\xe2\x9c\x8d',
	'x': '\xe2\x9d\x8c',
	'yarn': '\xf0\x9f\xa7\xb6',
	'yawning_face': '\xf0\x9f\xa5\xb1',
	'yellow_circle': '\xf0\x9f\x9f\xa1',
	'yellow_heart': '\xf0\x9f\x92\x9b',
	'yellow_square': '\xf0\x9f\x9f\xa8',
	'yemen': '\xf0\x9f\x87\xbe\xf0\x9f\x87\xaa',
	'yen': '\xf0\x9f\x92\xb4',
	'yin_yang': '\xe2\x98\xaf',
	'yo_yo': '\xf0\x9f\xaa\x80',
	'yum': '\xf0\x9f\x98\x8b',
	'zambia': '\xf0\x9f\x87\xbf\xf0\x9f\x87\xb2',
	'zany_face': '\xf0\x9f\xa4\xaa',
	'zap': '\xe2\x9a\xa1',
	'zebra': '\xf0\x9f\xa6\x93',
	'zero': '\x30\xe2\x83\xa3',
	'zimbabwe': '\xf0\x9f\x87\xbf\xf0\x9f\x87\xbc',
	'zipper_mouth_face': '\xf0\x9f\xa4\x90',
	'zombie': '\xf0\x9f\xa7\x9f',
	'zombie_man': '\xf0\x9f\xa7\x9f\xe2\x99\x82',
	'zombie_woman': '\xf0\x9f\xa7\x9f\xe2\x99\x80',
	'zzz': '\xf0\x9f\x92\xa4',
}
